`timescale 1 ns/100 ps
// Version: 2023.1 2023.1.0.6


module PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM(
       W_DATA,
       R_DATA,
       W_ADDR,
       R_ADDR,
       W_EN,
       R_EN,
       CLK,
       WBYTE_EN
    );
input  [39:0] W_DATA;
output [39:0] R_DATA;
input  [14:0] W_ADDR;
input  [14:0] R_ADDR;
input  W_EN;
input  R_EN;
input  CLK;
input  [3:0] WBYTE_EN;

    wire \R_DATA_TEMPR0[0] , \R_DATA_TEMPR1[0] , \R_DATA_TEMPR2[0] , 
        \R_DATA_TEMPR3[0] , \R_DATA_TEMPR4[0] , \R_DATA_TEMPR5[0] , 
        \R_DATA_TEMPR6[0] , \R_DATA_TEMPR7[0] , \R_DATA_TEMPR8[0] , 
        \R_DATA_TEMPR9[0] , \R_DATA_TEMPR10[0] , \R_DATA_TEMPR11[0] , 
        \R_DATA_TEMPR12[0] , \R_DATA_TEMPR13[0] , \R_DATA_TEMPR14[0] , 
        \R_DATA_TEMPR15[0] , \R_DATA_TEMPR16[0] , \R_DATA_TEMPR17[0] , 
        \R_DATA_TEMPR18[0] , \R_DATA_TEMPR19[0] , \R_DATA_TEMPR20[0] , 
        \R_DATA_TEMPR21[0] , \R_DATA_TEMPR22[0] , \R_DATA_TEMPR23[0] , 
        \R_DATA_TEMPR24[0] , \R_DATA_TEMPR25[0] , \R_DATA_TEMPR26[0] , 
        \R_DATA_TEMPR27[0] , \R_DATA_TEMPR28[0] , \R_DATA_TEMPR29[0] , 
        \R_DATA_TEMPR30[0] , \R_DATA_TEMPR31[0] , \R_DATA_TEMPR32[0] , 
        \R_DATA_TEMPR33[0] , \R_DATA_TEMPR34[0] , \R_DATA_TEMPR35[0] , 
        \R_DATA_TEMPR36[0] , \R_DATA_TEMPR37[0] , \R_DATA_TEMPR38[0] , 
        \R_DATA_TEMPR39[0] , \R_DATA_TEMPR40[0] , \R_DATA_TEMPR41[0] , 
        \R_DATA_TEMPR42[0] , \R_DATA_TEMPR43[0] , \R_DATA_TEMPR44[0] , 
        \R_DATA_TEMPR45[0] , \R_DATA_TEMPR46[0] , \R_DATA_TEMPR47[0] , 
        \R_DATA_TEMPR48[0] , \R_DATA_TEMPR49[0] , \R_DATA_TEMPR50[0] , 
        \R_DATA_TEMPR51[0] , \R_DATA_TEMPR52[0] , \R_DATA_TEMPR53[0] , 
        \R_DATA_TEMPR54[0] , \R_DATA_TEMPR55[0] , \R_DATA_TEMPR56[0] , 
        \R_DATA_TEMPR57[0] , \R_DATA_TEMPR58[0] , \R_DATA_TEMPR59[0] , 
        \R_DATA_TEMPR60[0] , \R_DATA_TEMPR61[0] , \R_DATA_TEMPR62[0] , 
        \R_DATA_TEMPR63[0] , \R_DATA_TEMPR0[1] , \R_DATA_TEMPR1[1] , 
        \R_DATA_TEMPR2[1] , \R_DATA_TEMPR3[1] , \R_DATA_TEMPR4[1] , 
        \R_DATA_TEMPR5[1] , \R_DATA_TEMPR6[1] , \R_DATA_TEMPR7[1] , 
        \R_DATA_TEMPR8[1] , \R_DATA_TEMPR9[1] , \R_DATA_TEMPR10[1] , 
        \R_DATA_TEMPR11[1] , \R_DATA_TEMPR12[1] , \R_DATA_TEMPR13[1] , 
        \R_DATA_TEMPR14[1] , \R_DATA_TEMPR15[1] , \R_DATA_TEMPR16[1] , 
        \R_DATA_TEMPR17[1] , \R_DATA_TEMPR18[1] , \R_DATA_TEMPR19[1] , 
        \R_DATA_TEMPR20[1] , \R_DATA_TEMPR21[1] , \R_DATA_TEMPR22[1] , 
        \R_DATA_TEMPR23[1] , \R_DATA_TEMPR24[1] , \R_DATA_TEMPR25[1] , 
        \R_DATA_TEMPR26[1] , \R_DATA_TEMPR27[1] , \R_DATA_TEMPR28[1] , 
        \R_DATA_TEMPR29[1] , \R_DATA_TEMPR30[1] , \R_DATA_TEMPR31[1] , 
        \R_DATA_TEMPR32[1] , \R_DATA_TEMPR33[1] , \R_DATA_TEMPR34[1] , 
        \R_DATA_TEMPR35[1] , \R_DATA_TEMPR36[1] , \R_DATA_TEMPR37[1] , 
        \R_DATA_TEMPR38[1] , \R_DATA_TEMPR39[1] , \R_DATA_TEMPR40[1] , 
        \R_DATA_TEMPR41[1] , \R_DATA_TEMPR42[1] , \R_DATA_TEMPR43[1] , 
        \R_DATA_TEMPR44[1] , \R_DATA_TEMPR45[1] , \R_DATA_TEMPR46[1] , 
        \R_DATA_TEMPR47[1] , \R_DATA_TEMPR48[1] , \R_DATA_TEMPR49[1] , 
        \R_DATA_TEMPR50[1] , \R_DATA_TEMPR51[1] , \R_DATA_TEMPR52[1] , 
        \R_DATA_TEMPR53[1] , \R_DATA_TEMPR54[1] , \R_DATA_TEMPR55[1] , 
        \R_DATA_TEMPR56[1] , \R_DATA_TEMPR57[1] , \R_DATA_TEMPR58[1] , 
        \R_DATA_TEMPR59[1] , \R_DATA_TEMPR60[1] , \R_DATA_TEMPR61[1] , 
        \R_DATA_TEMPR62[1] , \R_DATA_TEMPR63[1] , \R_DATA_TEMPR0[2] , 
        \R_DATA_TEMPR1[2] , \R_DATA_TEMPR2[2] , \R_DATA_TEMPR3[2] , 
        \R_DATA_TEMPR4[2] , \R_DATA_TEMPR5[2] , \R_DATA_TEMPR6[2] , 
        \R_DATA_TEMPR7[2] , \R_DATA_TEMPR8[2] , \R_DATA_TEMPR9[2] , 
        \R_DATA_TEMPR10[2] , \R_DATA_TEMPR11[2] , \R_DATA_TEMPR12[2] , 
        \R_DATA_TEMPR13[2] , \R_DATA_TEMPR14[2] , \R_DATA_TEMPR15[2] , 
        \R_DATA_TEMPR16[2] , \R_DATA_TEMPR17[2] , \R_DATA_TEMPR18[2] , 
        \R_DATA_TEMPR19[2] , \R_DATA_TEMPR20[2] , \R_DATA_TEMPR21[2] , 
        \R_DATA_TEMPR22[2] , \R_DATA_TEMPR23[2] , \R_DATA_TEMPR24[2] , 
        \R_DATA_TEMPR25[2] , \R_DATA_TEMPR26[2] , \R_DATA_TEMPR27[2] , 
        \R_DATA_TEMPR28[2] , \R_DATA_TEMPR29[2] , \R_DATA_TEMPR30[2] , 
        \R_DATA_TEMPR31[2] , \R_DATA_TEMPR32[2] , \R_DATA_TEMPR33[2] , 
        \R_DATA_TEMPR34[2] , \R_DATA_TEMPR35[2] , \R_DATA_TEMPR36[2] , 
        \R_DATA_TEMPR37[2] , \R_DATA_TEMPR38[2] , \R_DATA_TEMPR39[2] , 
        \R_DATA_TEMPR40[2] , \R_DATA_TEMPR41[2] , \R_DATA_TEMPR42[2] , 
        \R_DATA_TEMPR43[2] , \R_DATA_TEMPR44[2] , \R_DATA_TEMPR45[2] , 
        \R_DATA_TEMPR46[2] , \R_DATA_TEMPR47[2] , \R_DATA_TEMPR48[2] , 
        \R_DATA_TEMPR49[2] , \R_DATA_TEMPR50[2] , \R_DATA_TEMPR51[2] , 
        \R_DATA_TEMPR52[2] , \R_DATA_TEMPR53[2] , \R_DATA_TEMPR54[2] , 
        \R_DATA_TEMPR55[2] , \R_DATA_TEMPR56[2] , \R_DATA_TEMPR57[2] , 
        \R_DATA_TEMPR58[2] , \R_DATA_TEMPR59[2] , \R_DATA_TEMPR60[2] , 
        \R_DATA_TEMPR61[2] , \R_DATA_TEMPR62[2] , \R_DATA_TEMPR63[2] , 
        \R_DATA_TEMPR0[3] , \R_DATA_TEMPR1[3] , \R_DATA_TEMPR2[3] , 
        \R_DATA_TEMPR3[3] , \R_DATA_TEMPR4[3] , \R_DATA_TEMPR5[3] , 
        \R_DATA_TEMPR6[3] , \R_DATA_TEMPR7[3] , \R_DATA_TEMPR8[3] , 
        \R_DATA_TEMPR9[3] , \R_DATA_TEMPR10[3] , \R_DATA_TEMPR11[3] , 
        \R_DATA_TEMPR12[3] , \R_DATA_TEMPR13[3] , \R_DATA_TEMPR14[3] , 
        \R_DATA_TEMPR15[3] , \R_DATA_TEMPR16[3] , \R_DATA_TEMPR17[3] , 
        \R_DATA_TEMPR18[3] , \R_DATA_TEMPR19[3] , \R_DATA_TEMPR20[3] , 
        \R_DATA_TEMPR21[3] , \R_DATA_TEMPR22[3] , \R_DATA_TEMPR23[3] , 
        \R_DATA_TEMPR24[3] , \R_DATA_TEMPR25[3] , \R_DATA_TEMPR26[3] , 
        \R_DATA_TEMPR27[3] , \R_DATA_TEMPR28[3] , \R_DATA_TEMPR29[3] , 
        \R_DATA_TEMPR30[3] , \R_DATA_TEMPR31[3] , \R_DATA_TEMPR32[3] , 
        \R_DATA_TEMPR33[3] , \R_DATA_TEMPR34[3] , \R_DATA_TEMPR35[3] , 
        \R_DATA_TEMPR36[3] , \R_DATA_TEMPR37[3] , \R_DATA_TEMPR38[3] , 
        \R_DATA_TEMPR39[3] , \R_DATA_TEMPR40[3] , \R_DATA_TEMPR41[3] , 
        \R_DATA_TEMPR42[3] , \R_DATA_TEMPR43[3] , \R_DATA_TEMPR44[3] , 
        \R_DATA_TEMPR45[3] , \R_DATA_TEMPR46[3] , \R_DATA_TEMPR47[3] , 
        \R_DATA_TEMPR48[3] , \R_DATA_TEMPR49[3] , \R_DATA_TEMPR50[3] , 
        \R_DATA_TEMPR51[3] , \R_DATA_TEMPR52[3] , \R_DATA_TEMPR53[3] , 
        \R_DATA_TEMPR54[3] , \R_DATA_TEMPR55[3] , \R_DATA_TEMPR56[3] , 
        \R_DATA_TEMPR57[3] , \R_DATA_TEMPR58[3] , \R_DATA_TEMPR59[3] , 
        \R_DATA_TEMPR60[3] , \R_DATA_TEMPR61[3] , \R_DATA_TEMPR62[3] , 
        \R_DATA_TEMPR63[3] , \R_DATA_TEMPR0[4] , \R_DATA_TEMPR1[4] , 
        \R_DATA_TEMPR2[4] , \R_DATA_TEMPR3[4] , \R_DATA_TEMPR4[4] , 
        \R_DATA_TEMPR5[4] , \R_DATA_TEMPR6[4] , \R_DATA_TEMPR7[4] , 
        \R_DATA_TEMPR8[4] , \R_DATA_TEMPR9[4] , \R_DATA_TEMPR10[4] , 
        \R_DATA_TEMPR11[4] , \R_DATA_TEMPR12[4] , \R_DATA_TEMPR13[4] , 
        \R_DATA_TEMPR14[4] , \R_DATA_TEMPR15[4] , \R_DATA_TEMPR16[4] , 
        \R_DATA_TEMPR17[4] , \R_DATA_TEMPR18[4] , \R_DATA_TEMPR19[4] , 
        \R_DATA_TEMPR20[4] , \R_DATA_TEMPR21[4] , \R_DATA_TEMPR22[4] , 
        \R_DATA_TEMPR23[4] , \R_DATA_TEMPR24[4] , \R_DATA_TEMPR25[4] , 
        \R_DATA_TEMPR26[4] , \R_DATA_TEMPR27[4] , \R_DATA_TEMPR28[4] , 
        \R_DATA_TEMPR29[4] , \R_DATA_TEMPR30[4] , \R_DATA_TEMPR31[4] , 
        \R_DATA_TEMPR32[4] , \R_DATA_TEMPR33[4] , \R_DATA_TEMPR34[4] , 
        \R_DATA_TEMPR35[4] , \R_DATA_TEMPR36[4] , \R_DATA_TEMPR37[4] , 
        \R_DATA_TEMPR38[4] , \R_DATA_TEMPR39[4] , \R_DATA_TEMPR40[4] , 
        \R_DATA_TEMPR41[4] , \R_DATA_TEMPR42[4] , \R_DATA_TEMPR43[4] , 
        \R_DATA_TEMPR44[4] , \R_DATA_TEMPR45[4] , \R_DATA_TEMPR46[4] , 
        \R_DATA_TEMPR47[4] , \R_DATA_TEMPR48[4] , \R_DATA_TEMPR49[4] , 
        \R_DATA_TEMPR50[4] , \R_DATA_TEMPR51[4] , \R_DATA_TEMPR52[4] , 
        \R_DATA_TEMPR53[4] , \R_DATA_TEMPR54[4] , \R_DATA_TEMPR55[4] , 
        \R_DATA_TEMPR56[4] , \R_DATA_TEMPR57[4] , \R_DATA_TEMPR58[4] , 
        \R_DATA_TEMPR59[4] , \R_DATA_TEMPR60[4] , \R_DATA_TEMPR61[4] , 
        \R_DATA_TEMPR62[4] , \R_DATA_TEMPR63[4] , \R_DATA_TEMPR0[5] , 
        \R_DATA_TEMPR1[5] , \R_DATA_TEMPR2[5] , \R_DATA_TEMPR3[5] , 
        \R_DATA_TEMPR4[5] , \R_DATA_TEMPR5[5] , \R_DATA_TEMPR6[5] , 
        \R_DATA_TEMPR7[5] , \R_DATA_TEMPR8[5] , \R_DATA_TEMPR9[5] , 
        \R_DATA_TEMPR10[5] , \R_DATA_TEMPR11[5] , \R_DATA_TEMPR12[5] , 
        \R_DATA_TEMPR13[5] , \R_DATA_TEMPR14[5] , \R_DATA_TEMPR15[5] , 
        \R_DATA_TEMPR16[5] , \R_DATA_TEMPR17[5] , \R_DATA_TEMPR18[5] , 
        \R_DATA_TEMPR19[5] , \R_DATA_TEMPR20[5] , \R_DATA_TEMPR21[5] , 
        \R_DATA_TEMPR22[5] , \R_DATA_TEMPR23[5] , \R_DATA_TEMPR24[5] , 
        \R_DATA_TEMPR25[5] , \R_DATA_TEMPR26[5] , \R_DATA_TEMPR27[5] , 
        \R_DATA_TEMPR28[5] , \R_DATA_TEMPR29[5] , \R_DATA_TEMPR30[5] , 
        \R_DATA_TEMPR31[5] , \R_DATA_TEMPR32[5] , \R_DATA_TEMPR33[5] , 
        \R_DATA_TEMPR34[5] , \R_DATA_TEMPR35[5] , \R_DATA_TEMPR36[5] , 
        \R_DATA_TEMPR37[5] , \R_DATA_TEMPR38[5] , \R_DATA_TEMPR39[5] , 
        \R_DATA_TEMPR40[5] , \R_DATA_TEMPR41[5] , \R_DATA_TEMPR42[5] , 
        \R_DATA_TEMPR43[5] , \R_DATA_TEMPR44[5] , \R_DATA_TEMPR45[5] , 
        \R_DATA_TEMPR46[5] , \R_DATA_TEMPR47[5] , \R_DATA_TEMPR48[5] , 
        \R_DATA_TEMPR49[5] , \R_DATA_TEMPR50[5] , \R_DATA_TEMPR51[5] , 
        \R_DATA_TEMPR52[5] , \R_DATA_TEMPR53[5] , \R_DATA_TEMPR54[5] , 
        \R_DATA_TEMPR55[5] , \R_DATA_TEMPR56[5] , \R_DATA_TEMPR57[5] , 
        \R_DATA_TEMPR58[5] , \R_DATA_TEMPR59[5] , \R_DATA_TEMPR60[5] , 
        \R_DATA_TEMPR61[5] , \R_DATA_TEMPR62[5] , \R_DATA_TEMPR63[5] , 
        \R_DATA_TEMPR0[6] , \R_DATA_TEMPR1[6] , \R_DATA_TEMPR2[6] , 
        \R_DATA_TEMPR3[6] , \R_DATA_TEMPR4[6] , \R_DATA_TEMPR5[6] , 
        \R_DATA_TEMPR6[6] , \R_DATA_TEMPR7[6] , \R_DATA_TEMPR8[6] , 
        \R_DATA_TEMPR9[6] , \R_DATA_TEMPR10[6] , \R_DATA_TEMPR11[6] , 
        \R_DATA_TEMPR12[6] , \R_DATA_TEMPR13[6] , \R_DATA_TEMPR14[6] , 
        \R_DATA_TEMPR15[6] , \R_DATA_TEMPR16[6] , \R_DATA_TEMPR17[6] , 
        \R_DATA_TEMPR18[6] , \R_DATA_TEMPR19[6] , \R_DATA_TEMPR20[6] , 
        \R_DATA_TEMPR21[6] , \R_DATA_TEMPR22[6] , \R_DATA_TEMPR23[6] , 
        \R_DATA_TEMPR24[6] , \R_DATA_TEMPR25[6] , \R_DATA_TEMPR26[6] , 
        \R_DATA_TEMPR27[6] , \R_DATA_TEMPR28[6] , \R_DATA_TEMPR29[6] , 
        \R_DATA_TEMPR30[6] , \R_DATA_TEMPR31[6] , \R_DATA_TEMPR32[6] , 
        \R_DATA_TEMPR33[6] , \R_DATA_TEMPR34[6] , \R_DATA_TEMPR35[6] , 
        \R_DATA_TEMPR36[6] , \R_DATA_TEMPR37[6] , \R_DATA_TEMPR38[6] , 
        \R_DATA_TEMPR39[6] , \R_DATA_TEMPR40[6] , \R_DATA_TEMPR41[6] , 
        \R_DATA_TEMPR42[6] , \R_DATA_TEMPR43[6] , \R_DATA_TEMPR44[6] , 
        \R_DATA_TEMPR45[6] , \R_DATA_TEMPR46[6] , \R_DATA_TEMPR47[6] , 
        \R_DATA_TEMPR48[6] , \R_DATA_TEMPR49[6] , \R_DATA_TEMPR50[6] , 
        \R_DATA_TEMPR51[6] , \R_DATA_TEMPR52[6] , \R_DATA_TEMPR53[6] , 
        \R_DATA_TEMPR54[6] , \R_DATA_TEMPR55[6] , \R_DATA_TEMPR56[6] , 
        \R_DATA_TEMPR57[6] , \R_DATA_TEMPR58[6] , \R_DATA_TEMPR59[6] , 
        \R_DATA_TEMPR60[6] , \R_DATA_TEMPR61[6] , \R_DATA_TEMPR62[6] , 
        \R_DATA_TEMPR63[6] , \R_DATA_TEMPR0[7] , \R_DATA_TEMPR1[7] , 
        \R_DATA_TEMPR2[7] , \R_DATA_TEMPR3[7] , \R_DATA_TEMPR4[7] , 
        \R_DATA_TEMPR5[7] , \R_DATA_TEMPR6[7] , \R_DATA_TEMPR7[7] , 
        \R_DATA_TEMPR8[7] , \R_DATA_TEMPR9[7] , \R_DATA_TEMPR10[7] , 
        \R_DATA_TEMPR11[7] , \R_DATA_TEMPR12[7] , \R_DATA_TEMPR13[7] , 
        \R_DATA_TEMPR14[7] , \R_DATA_TEMPR15[7] , \R_DATA_TEMPR16[7] , 
        \R_DATA_TEMPR17[7] , \R_DATA_TEMPR18[7] , \R_DATA_TEMPR19[7] , 
        \R_DATA_TEMPR20[7] , \R_DATA_TEMPR21[7] , \R_DATA_TEMPR22[7] , 
        \R_DATA_TEMPR23[7] , \R_DATA_TEMPR24[7] , \R_DATA_TEMPR25[7] , 
        \R_DATA_TEMPR26[7] , \R_DATA_TEMPR27[7] , \R_DATA_TEMPR28[7] , 
        \R_DATA_TEMPR29[7] , \R_DATA_TEMPR30[7] , \R_DATA_TEMPR31[7] , 
        \R_DATA_TEMPR32[7] , \R_DATA_TEMPR33[7] , \R_DATA_TEMPR34[7] , 
        \R_DATA_TEMPR35[7] , \R_DATA_TEMPR36[7] , \R_DATA_TEMPR37[7] , 
        \R_DATA_TEMPR38[7] , \R_DATA_TEMPR39[7] , \R_DATA_TEMPR40[7] , 
        \R_DATA_TEMPR41[7] , \R_DATA_TEMPR42[7] , \R_DATA_TEMPR43[7] , 
        \R_DATA_TEMPR44[7] , \R_DATA_TEMPR45[7] , \R_DATA_TEMPR46[7] , 
        \R_DATA_TEMPR47[7] , \R_DATA_TEMPR48[7] , \R_DATA_TEMPR49[7] , 
        \R_DATA_TEMPR50[7] , \R_DATA_TEMPR51[7] , \R_DATA_TEMPR52[7] , 
        \R_DATA_TEMPR53[7] , \R_DATA_TEMPR54[7] , \R_DATA_TEMPR55[7] , 
        \R_DATA_TEMPR56[7] , \R_DATA_TEMPR57[7] , \R_DATA_TEMPR58[7] , 
        \R_DATA_TEMPR59[7] , \R_DATA_TEMPR60[7] , \R_DATA_TEMPR61[7] , 
        \R_DATA_TEMPR62[7] , \R_DATA_TEMPR63[7] , \R_DATA_TEMPR0[8] , 
        \R_DATA_TEMPR1[8] , \R_DATA_TEMPR2[8] , \R_DATA_TEMPR3[8] , 
        \R_DATA_TEMPR4[8] , \R_DATA_TEMPR5[8] , \R_DATA_TEMPR6[8] , 
        \R_DATA_TEMPR7[8] , \R_DATA_TEMPR8[8] , \R_DATA_TEMPR9[8] , 
        \R_DATA_TEMPR10[8] , \R_DATA_TEMPR11[8] , \R_DATA_TEMPR12[8] , 
        \R_DATA_TEMPR13[8] , \R_DATA_TEMPR14[8] , \R_DATA_TEMPR15[8] , 
        \R_DATA_TEMPR16[8] , \R_DATA_TEMPR17[8] , \R_DATA_TEMPR18[8] , 
        \R_DATA_TEMPR19[8] , \R_DATA_TEMPR20[8] , \R_DATA_TEMPR21[8] , 
        \R_DATA_TEMPR22[8] , \R_DATA_TEMPR23[8] , \R_DATA_TEMPR24[8] , 
        \R_DATA_TEMPR25[8] , \R_DATA_TEMPR26[8] , \R_DATA_TEMPR27[8] , 
        \R_DATA_TEMPR28[8] , \R_DATA_TEMPR29[8] , \R_DATA_TEMPR30[8] , 
        \R_DATA_TEMPR31[8] , \R_DATA_TEMPR32[8] , \R_DATA_TEMPR33[8] , 
        \R_DATA_TEMPR34[8] , \R_DATA_TEMPR35[8] , \R_DATA_TEMPR36[8] , 
        \R_DATA_TEMPR37[8] , \R_DATA_TEMPR38[8] , \R_DATA_TEMPR39[8] , 
        \R_DATA_TEMPR40[8] , \R_DATA_TEMPR41[8] , \R_DATA_TEMPR42[8] , 
        \R_DATA_TEMPR43[8] , \R_DATA_TEMPR44[8] , \R_DATA_TEMPR45[8] , 
        \R_DATA_TEMPR46[8] , \R_DATA_TEMPR47[8] , \R_DATA_TEMPR48[8] , 
        \R_DATA_TEMPR49[8] , \R_DATA_TEMPR50[8] , \R_DATA_TEMPR51[8] , 
        \R_DATA_TEMPR52[8] , \R_DATA_TEMPR53[8] , \R_DATA_TEMPR54[8] , 
        \R_DATA_TEMPR55[8] , \R_DATA_TEMPR56[8] , \R_DATA_TEMPR57[8] , 
        \R_DATA_TEMPR58[8] , \R_DATA_TEMPR59[8] , \R_DATA_TEMPR60[8] , 
        \R_DATA_TEMPR61[8] , \R_DATA_TEMPR62[8] , \R_DATA_TEMPR63[8] , 
        \R_DATA_TEMPR0[9] , \R_DATA_TEMPR1[9] , \R_DATA_TEMPR2[9] , 
        \R_DATA_TEMPR3[9] , \R_DATA_TEMPR4[9] , \R_DATA_TEMPR5[9] , 
        \R_DATA_TEMPR6[9] , \R_DATA_TEMPR7[9] , \R_DATA_TEMPR8[9] , 
        \R_DATA_TEMPR9[9] , \R_DATA_TEMPR10[9] , \R_DATA_TEMPR11[9] , 
        \R_DATA_TEMPR12[9] , \R_DATA_TEMPR13[9] , \R_DATA_TEMPR14[9] , 
        \R_DATA_TEMPR15[9] , \R_DATA_TEMPR16[9] , \R_DATA_TEMPR17[9] , 
        \R_DATA_TEMPR18[9] , \R_DATA_TEMPR19[9] , \R_DATA_TEMPR20[9] , 
        \R_DATA_TEMPR21[9] , \R_DATA_TEMPR22[9] , \R_DATA_TEMPR23[9] , 
        \R_DATA_TEMPR24[9] , \R_DATA_TEMPR25[9] , \R_DATA_TEMPR26[9] , 
        \R_DATA_TEMPR27[9] , \R_DATA_TEMPR28[9] , \R_DATA_TEMPR29[9] , 
        \R_DATA_TEMPR30[9] , \R_DATA_TEMPR31[9] , \R_DATA_TEMPR32[9] , 
        \R_DATA_TEMPR33[9] , \R_DATA_TEMPR34[9] , \R_DATA_TEMPR35[9] , 
        \R_DATA_TEMPR36[9] , \R_DATA_TEMPR37[9] , \R_DATA_TEMPR38[9] , 
        \R_DATA_TEMPR39[9] , \R_DATA_TEMPR40[9] , \R_DATA_TEMPR41[9] , 
        \R_DATA_TEMPR42[9] , \R_DATA_TEMPR43[9] , \R_DATA_TEMPR44[9] , 
        \R_DATA_TEMPR45[9] , \R_DATA_TEMPR46[9] , \R_DATA_TEMPR47[9] , 
        \R_DATA_TEMPR48[9] , \R_DATA_TEMPR49[9] , \R_DATA_TEMPR50[9] , 
        \R_DATA_TEMPR51[9] , \R_DATA_TEMPR52[9] , \R_DATA_TEMPR53[9] , 
        \R_DATA_TEMPR54[9] , \R_DATA_TEMPR55[9] , \R_DATA_TEMPR56[9] , 
        \R_DATA_TEMPR57[9] , \R_DATA_TEMPR58[9] , \R_DATA_TEMPR59[9] , 
        \R_DATA_TEMPR60[9] , \R_DATA_TEMPR61[9] , \R_DATA_TEMPR62[9] , 
        \R_DATA_TEMPR63[9] , \R_DATA_TEMPR0[10] , \R_DATA_TEMPR1[10] , 
        \R_DATA_TEMPR2[10] , \R_DATA_TEMPR3[10] , \R_DATA_TEMPR4[10] , 
        \R_DATA_TEMPR5[10] , \R_DATA_TEMPR6[10] , \R_DATA_TEMPR7[10] , 
        \R_DATA_TEMPR8[10] , \R_DATA_TEMPR9[10] , \R_DATA_TEMPR10[10] , 
        \R_DATA_TEMPR11[10] , \R_DATA_TEMPR12[10] , 
        \R_DATA_TEMPR13[10] , \R_DATA_TEMPR14[10] , 
        \R_DATA_TEMPR15[10] , \R_DATA_TEMPR16[10] , 
        \R_DATA_TEMPR17[10] , \R_DATA_TEMPR18[10] , 
        \R_DATA_TEMPR19[10] , \R_DATA_TEMPR20[10] , 
        \R_DATA_TEMPR21[10] , \R_DATA_TEMPR22[10] , 
        \R_DATA_TEMPR23[10] , \R_DATA_TEMPR24[10] , 
        \R_DATA_TEMPR25[10] , \R_DATA_TEMPR26[10] , 
        \R_DATA_TEMPR27[10] , \R_DATA_TEMPR28[10] , 
        \R_DATA_TEMPR29[10] , \R_DATA_TEMPR30[10] , 
        \R_DATA_TEMPR31[10] , \R_DATA_TEMPR32[10] , 
        \R_DATA_TEMPR33[10] , \R_DATA_TEMPR34[10] , 
        \R_DATA_TEMPR35[10] , \R_DATA_TEMPR36[10] , 
        \R_DATA_TEMPR37[10] , \R_DATA_TEMPR38[10] , 
        \R_DATA_TEMPR39[10] , \R_DATA_TEMPR40[10] , 
        \R_DATA_TEMPR41[10] , \R_DATA_TEMPR42[10] , 
        \R_DATA_TEMPR43[10] , \R_DATA_TEMPR44[10] , 
        \R_DATA_TEMPR45[10] , \R_DATA_TEMPR46[10] , 
        \R_DATA_TEMPR47[10] , \R_DATA_TEMPR48[10] , 
        \R_DATA_TEMPR49[10] , \R_DATA_TEMPR50[10] , 
        \R_DATA_TEMPR51[10] , \R_DATA_TEMPR52[10] , 
        \R_DATA_TEMPR53[10] , \R_DATA_TEMPR54[10] , 
        \R_DATA_TEMPR55[10] , \R_DATA_TEMPR56[10] , 
        \R_DATA_TEMPR57[10] , \R_DATA_TEMPR58[10] , 
        \R_DATA_TEMPR59[10] , \R_DATA_TEMPR60[10] , 
        \R_DATA_TEMPR61[10] , \R_DATA_TEMPR62[10] , 
        \R_DATA_TEMPR63[10] , \R_DATA_TEMPR0[11] , \R_DATA_TEMPR1[11] , 
        \R_DATA_TEMPR2[11] , \R_DATA_TEMPR3[11] , \R_DATA_TEMPR4[11] , 
        \R_DATA_TEMPR5[11] , \R_DATA_TEMPR6[11] , \R_DATA_TEMPR7[11] , 
        \R_DATA_TEMPR8[11] , \R_DATA_TEMPR9[11] , \R_DATA_TEMPR10[11] , 
        \R_DATA_TEMPR11[11] , \R_DATA_TEMPR12[11] , 
        \R_DATA_TEMPR13[11] , \R_DATA_TEMPR14[11] , 
        \R_DATA_TEMPR15[11] , \R_DATA_TEMPR16[11] , 
        \R_DATA_TEMPR17[11] , \R_DATA_TEMPR18[11] , 
        \R_DATA_TEMPR19[11] , \R_DATA_TEMPR20[11] , 
        \R_DATA_TEMPR21[11] , \R_DATA_TEMPR22[11] , 
        \R_DATA_TEMPR23[11] , \R_DATA_TEMPR24[11] , 
        \R_DATA_TEMPR25[11] , \R_DATA_TEMPR26[11] , 
        \R_DATA_TEMPR27[11] , \R_DATA_TEMPR28[11] , 
        \R_DATA_TEMPR29[11] , \R_DATA_TEMPR30[11] , 
        \R_DATA_TEMPR31[11] , \R_DATA_TEMPR32[11] , 
        \R_DATA_TEMPR33[11] , \R_DATA_TEMPR34[11] , 
        \R_DATA_TEMPR35[11] , \R_DATA_TEMPR36[11] , 
        \R_DATA_TEMPR37[11] , \R_DATA_TEMPR38[11] , 
        \R_DATA_TEMPR39[11] , \R_DATA_TEMPR40[11] , 
        \R_DATA_TEMPR41[11] , \R_DATA_TEMPR42[11] , 
        \R_DATA_TEMPR43[11] , \R_DATA_TEMPR44[11] , 
        \R_DATA_TEMPR45[11] , \R_DATA_TEMPR46[11] , 
        \R_DATA_TEMPR47[11] , \R_DATA_TEMPR48[11] , 
        \R_DATA_TEMPR49[11] , \R_DATA_TEMPR50[11] , 
        \R_DATA_TEMPR51[11] , \R_DATA_TEMPR52[11] , 
        \R_DATA_TEMPR53[11] , \R_DATA_TEMPR54[11] , 
        \R_DATA_TEMPR55[11] , \R_DATA_TEMPR56[11] , 
        \R_DATA_TEMPR57[11] , \R_DATA_TEMPR58[11] , 
        \R_DATA_TEMPR59[11] , \R_DATA_TEMPR60[11] , 
        \R_DATA_TEMPR61[11] , \R_DATA_TEMPR62[11] , 
        \R_DATA_TEMPR63[11] , \R_DATA_TEMPR0[12] , \R_DATA_TEMPR1[12] , 
        \R_DATA_TEMPR2[12] , \R_DATA_TEMPR3[12] , \R_DATA_TEMPR4[12] , 
        \R_DATA_TEMPR5[12] , \R_DATA_TEMPR6[12] , \R_DATA_TEMPR7[12] , 
        \R_DATA_TEMPR8[12] , \R_DATA_TEMPR9[12] , \R_DATA_TEMPR10[12] , 
        \R_DATA_TEMPR11[12] , \R_DATA_TEMPR12[12] , 
        \R_DATA_TEMPR13[12] , \R_DATA_TEMPR14[12] , 
        \R_DATA_TEMPR15[12] , \R_DATA_TEMPR16[12] , 
        \R_DATA_TEMPR17[12] , \R_DATA_TEMPR18[12] , 
        \R_DATA_TEMPR19[12] , \R_DATA_TEMPR20[12] , 
        \R_DATA_TEMPR21[12] , \R_DATA_TEMPR22[12] , 
        \R_DATA_TEMPR23[12] , \R_DATA_TEMPR24[12] , 
        \R_DATA_TEMPR25[12] , \R_DATA_TEMPR26[12] , 
        \R_DATA_TEMPR27[12] , \R_DATA_TEMPR28[12] , 
        \R_DATA_TEMPR29[12] , \R_DATA_TEMPR30[12] , 
        \R_DATA_TEMPR31[12] , \R_DATA_TEMPR32[12] , 
        \R_DATA_TEMPR33[12] , \R_DATA_TEMPR34[12] , 
        \R_DATA_TEMPR35[12] , \R_DATA_TEMPR36[12] , 
        \R_DATA_TEMPR37[12] , \R_DATA_TEMPR38[12] , 
        \R_DATA_TEMPR39[12] , \R_DATA_TEMPR40[12] , 
        \R_DATA_TEMPR41[12] , \R_DATA_TEMPR42[12] , 
        \R_DATA_TEMPR43[12] , \R_DATA_TEMPR44[12] , 
        \R_DATA_TEMPR45[12] , \R_DATA_TEMPR46[12] , 
        \R_DATA_TEMPR47[12] , \R_DATA_TEMPR48[12] , 
        \R_DATA_TEMPR49[12] , \R_DATA_TEMPR50[12] , 
        \R_DATA_TEMPR51[12] , \R_DATA_TEMPR52[12] , 
        \R_DATA_TEMPR53[12] , \R_DATA_TEMPR54[12] , 
        \R_DATA_TEMPR55[12] , \R_DATA_TEMPR56[12] , 
        \R_DATA_TEMPR57[12] , \R_DATA_TEMPR58[12] , 
        \R_DATA_TEMPR59[12] , \R_DATA_TEMPR60[12] , 
        \R_DATA_TEMPR61[12] , \R_DATA_TEMPR62[12] , 
        \R_DATA_TEMPR63[12] , \R_DATA_TEMPR0[13] , \R_DATA_TEMPR1[13] , 
        \R_DATA_TEMPR2[13] , \R_DATA_TEMPR3[13] , \R_DATA_TEMPR4[13] , 
        \R_DATA_TEMPR5[13] , \R_DATA_TEMPR6[13] , \R_DATA_TEMPR7[13] , 
        \R_DATA_TEMPR8[13] , \R_DATA_TEMPR9[13] , \R_DATA_TEMPR10[13] , 
        \R_DATA_TEMPR11[13] , \R_DATA_TEMPR12[13] , 
        \R_DATA_TEMPR13[13] , \R_DATA_TEMPR14[13] , 
        \R_DATA_TEMPR15[13] , \R_DATA_TEMPR16[13] , 
        \R_DATA_TEMPR17[13] , \R_DATA_TEMPR18[13] , 
        \R_DATA_TEMPR19[13] , \R_DATA_TEMPR20[13] , 
        \R_DATA_TEMPR21[13] , \R_DATA_TEMPR22[13] , 
        \R_DATA_TEMPR23[13] , \R_DATA_TEMPR24[13] , 
        \R_DATA_TEMPR25[13] , \R_DATA_TEMPR26[13] , 
        \R_DATA_TEMPR27[13] , \R_DATA_TEMPR28[13] , 
        \R_DATA_TEMPR29[13] , \R_DATA_TEMPR30[13] , 
        \R_DATA_TEMPR31[13] , \R_DATA_TEMPR32[13] , 
        \R_DATA_TEMPR33[13] , \R_DATA_TEMPR34[13] , 
        \R_DATA_TEMPR35[13] , \R_DATA_TEMPR36[13] , 
        \R_DATA_TEMPR37[13] , \R_DATA_TEMPR38[13] , 
        \R_DATA_TEMPR39[13] , \R_DATA_TEMPR40[13] , 
        \R_DATA_TEMPR41[13] , \R_DATA_TEMPR42[13] , 
        \R_DATA_TEMPR43[13] , \R_DATA_TEMPR44[13] , 
        \R_DATA_TEMPR45[13] , \R_DATA_TEMPR46[13] , 
        \R_DATA_TEMPR47[13] , \R_DATA_TEMPR48[13] , 
        \R_DATA_TEMPR49[13] , \R_DATA_TEMPR50[13] , 
        \R_DATA_TEMPR51[13] , \R_DATA_TEMPR52[13] , 
        \R_DATA_TEMPR53[13] , \R_DATA_TEMPR54[13] , 
        \R_DATA_TEMPR55[13] , \R_DATA_TEMPR56[13] , 
        \R_DATA_TEMPR57[13] , \R_DATA_TEMPR58[13] , 
        \R_DATA_TEMPR59[13] , \R_DATA_TEMPR60[13] , 
        \R_DATA_TEMPR61[13] , \R_DATA_TEMPR62[13] , 
        \R_DATA_TEMPR63[13] , \R_DATA_TEMPR0[14] , \R_DATA_TEMPR1[14] , 
        \R_DATA_TEMPR2[14] , \R_DATA_TEMPR3[14] , \R_DATA_TEMPR4[14] , 
        \R_DATA_TEMPR5[14] , \R_DATA_TEMPR6[14] , \R_DATA_TEMPR7[14] , 
        \R_DATA_TEMPR8[14] , \R_DATA_TEMPR9[14] , \R_DATA_TEMPR10[14] , 
        \R_DATA_TEMPR11[14] , \R_DATA_TEMPR12[14] , 
        \R_DATA_TEMPR13[14] , \R_DATA_TEMPR14[14] , 
        \R_DATA_TEMPR15[14] , \R_DATA_TEMPR16[14] , 
        \R_DATA_TEMPR17[14] , \R_DATA_TEMPR18[14] , 
        \R_DATA_TEMPR19[14] , \R_DATA_TEMPR20[14] , 
        \R_DATA_TEMPR21[14] , \R_DATA_TEMPR22[14] , 
        \R_DATA_TEMPR23[14] , \R_DATA_TEMPR24[14] , 
        \R_DATA_TEMPR25[14] , \R_DATA_TEMPR26[14] , 
        \R_DATA_TEMPR27[14] , \R_DATA_TEMPR28[14] , 
        \R_DATA_TEMPR29[14] , \R_DATA_TEMPR30[14] , 
        \R_DATA_TEMPR31[14] , \R_DATA_TEMPR32[14] , 
        \R_DATA_TEMPR33[14] , \R_DATA_TEMPR34[14] , 
        \R_DATA_TEMPR35[14] , \R_DATA_TEMPR36[14] , 
        \R_DATA_TEMPR37[14] , \R_DATA_TEMPR38[14] , 
        \R_DATA_TEMPR39[14] , \R_DATA_TEMPR40[14] , 
        \R_DATA_TEMPR41[14] , \R_DATA_TEMPR42[14] , 
        \R_DATA_TEMPR43[14] , \R_DATA_TEMPR44[14] , 
        \R_DATA_TEMPR45[14] , \R_DATA_TEMPR46[14] , 
        \R_DATA_TEMPR47[14] , \R_DATA_TEMPR48[14] , 
        \R_DATA_TEMPR49[14] , \R_DATA_TEMPR50[14] , 
        \R_DATA_TEMPR51[14] , \R_DATA_TEMPR52[14] , 
        \R_DATA_TEMPR53[14] , \R_DATA_TEMPR54[14] , 
        \R_DATA_TEMPR55[14] , \R_DATA_TEMPR56[14] , 
        \R_DATA_TEMPR57[14] , \R_DATA_TEMPR58[14] , 
        \R_DATA_TEMPR59[14] , \R_DATA_TEMPR60[14] , 
        \R_DATA_TEMPR61[14] , \R_DATA_TEMPR62[14] , 
        \R_DATA_TEMPR63[14] , \R_DATA_TEMPR0[15] , \R_DATA_TEMPR1[15] , 
        \R_DATA_TEMPR2[15] , \R_DATA_TEMPR3[15] , \R_DATA_TEMPR4[15] , 
        \R_DATA_TEMPR5[15] , \R_DATA_TEMPR6[15] , \R_DATA_TEMPR7[15] , 
        \R_DATA_TEMPR8[15] , \R_DATA_TEMPR9[15] , \R_DATA_TEMPR10[15] , 
        \R_DATA_TEMPR11[15] , \R_DATA_TEMPR12[15] , 
        \R_DATA_TEMPR13[15] , \R_DATA_TEMPR14[15] , 
        \R_DATA_TEMPR15[15] , \R_DATA_TEMPR16[15] , 
        \R_DATA_TEMPR17[15] , \R_DATA_TEMPR18[15] , 
        \R_DATA_TEMPR19[15] , \R_DATA_TEMPR20[15] , 
        \R_DATA_TEMPR21[15] , \R_DATA_TEMPR22[15] , 
        \R_DATA_TEMPR23[15] , \R_DATA_TEMPR24[15] , 
        \R_DATA_TEMPR25[15] , \R_DATA_TEMPR26[15] , 
        \R_DATA_TEMPR27[15] , \R_DATA_TEMPR28[15] , 
        \R_DATA_TEMPR29[15] , \R_DATA_TEMPR30[15] , 
        \R_DATA_TEMPR31[15] , \R_DATA_TEMPR32[15] , 
        \R_DATA_TEMPR33[15] , \R_DATA_TEMPR34[15] , 
        \R_DATA_TEMPR35[15] , \R_DATA_TEMPR36[15] , 
        \R_DATA_TEMPR37[15] , \R_DATA_TEMPR38[15] , 
        \R_DATA_TEMPR39[15] , \R_DATA_TEMPR40[15] , 
        \R_DATA_TEMPR41[15] , \R_DATA_TEMPR42[15] , 
        \R_DATA_TEMPR43[15] , \R_DATA_TEMPR44[15] , 
        \R_DATA_TEMPR45[15] , \R_DATA_TEMPR46[15] , 
        \R_DATA_TEMPR47[15] , \R_DATA_TEMPR48[15] , 
        \R_DATA_TEMPR49[15] , \R_DATA_TEMPR50[15] , 
        \R_DATA_TEMPR51[15] , \R_DATA_TEMPR52[15] , 
        \R_DATA_TEMPR53[15] , \R_DATA_TEMPR54[15] , 
        \R_DATA_TEMPR55[15] , \R_DATA_TEMPR56[15] , 
        \R_DATA_TEMPR57[15] , \R_DATA_TEMPR58[15] , 
        \R_DATA_TEMPR59[15] , \R_DATA_TEMPR60[15] , 
        \R_DATA_TEMPR61[15] , \R_DATA_TEMPR62[15] , 
        \R_DATA_TEMPR63[15] , \R_DATA_TEMPR0[16] , \R_DATA_TEMPR1[16] , 
        \R_DATA_TEMPR2[16] , \R_DATA_TEMPR3[16] , \R_DATA_TEMPR4[16] , 
        \R_DATA_TEMPR5[16] , \R_DATA_TEMPR6[16] , \R_DATA_TEMPR7[16] , 
        \R_DATA_TEMPR8[16] , \R_DATA_TEMPR9[16] , \R_DATA_TEMPR10[16] , 
        \R_DATA_TEMPR11[16] , \R_DATA_TEMPR12[16] , 
        \R_DATA_TEMPR13[16] , \R_DATA_TEMPR14[16] , 
        \R_DATA_TEMPR15[16] , \R_DATA_TEMPR16[16] , 
        \R_DATA_TEMPR17[16] , \R_DATA_TEMPR18[16] , 
        \R_DATA_TEMPR19[16] , \R_DATA_TEMPR20[16] , 
        \R_DATA_TEMPR21[16] , \R_DATA_TEMPR22[16] , 
        \R_DATA_TEMPR23[16] , \R_DATA_TEMPR24[16] , 
        \R_DATA_TEMPR25[16] , \R_DATA_TEMPR26[16] , 
        \R_DATA_TEMPR27[16] , \R_DATA_TEMPR28[16] , 
        \R_DATA_TEMPR29[16] , \R_DATA_TEMPR30[16] , 
        \R_DATA_TEMPR31[16] , \R_DATA_TEMPR32[16] , 
        \R_DATA_TEMPR33[16] , \R_DATA_TEMPR34[16] , 
        \R_DATA_TEMPR35[16] , \R_DATA_TEMPR36[16] , 
        \R_DATA_TEMPR37[16] , \R_DATA_TEMPR38[16] , 
        \R_DATA_TEMPR39[16] , \R_DATA_TEMPR40[16] , 
        \R_DATA_TEMPR41[16] , \R_DATA_TEMPR42[16] , 
        \R_DATA_TEMPR43[16] , \R_DATA_TEMPR44[16] , 
        \R_DATA_TEMPR45[16] , \R_DATA_TEMPR46[16] , 
        \R_DATA_TEMPR47[16] , \R_DATA_TEMPR48[16] , 
        \R_DATA_TEMPR49[16] , \R_DATA_TEMPR50[16] , 
        \R_DATA_TEMPR51[16] , \R_DATA_TEMPR52[16] , 
        \R_DATA_TEMPR53[16] , \R_DATA_TEMPR54[16] , 
        \R_DATA_TEMPR55[16] , \R_DATA_TEMPR56[16] , 
        \R_DATA_TEMPR57[16] , \R_DATA_TEMPR58[16] , 
        \R_DATA_TEMPR59[16] , \R_DATA_TEMPR60[16] , 
        \R_DATA_TEMPR61[16] , \R_DATA_TEMPR62[16] , 
        \R_DATA_TEMPR63[16] , \R_DATA_TEMPR0[17] , \R_DATA_TEMPR1[17] , 
        \R_DATA_TEMPR2[17] , \R_DATA_TEMPR3[17] , \R_DATA_TEMPR4[17] , 
        \R_DATA_TEMPR5[17] , \R_DATA_TEMPR6[17] , \R_DATA_TEMPR7[17] , 
        \R_DATA_TEMPR8[17] , \R_DATA_TEMPR9[17] , \R_DATA_TEMPR10[17] , 
        \R_DATA_TEMPR11[17] , \R_DATA_TEMPR12[17] , 
        \R_DATA_TEMPR13[17] , \R_DATA_TEMPR14[17] , 
        \R_DATA_TEMPR15[17] , \R_DATA_TEMPR16[17] , 
        \R_DATA_TEMPR17[17] , \R_DATA_TEMPR18[17] , 
        \R_DATA_TEMPR19[17] , \R_DATA_TEMPR20[17] , 
        \R_DATA_TEMPR21[17] , \R_DATA_TEMPR22[17] , 
        \R_DATA_TEMPR23[17] , \R_DATA_TEMPR24[17] , 
        \R_DATA_TEMPR25[17] , \R_DATA_TEMPR26[17] , 
        \R_DATA_TEMPR27[17] , \R_DATA_TEMPR28[17] , 
        \R_DATA_TEMPR29[17] , \R_DATA_TEMPR30[17] , 
        \R_DATA_TEMPR31[17] , \R_DATA_TEMPR32[17] , 
        \R_DATA_TEMPR33[17] , \R_DATA_TEMPR34[17] , 
        \R_DATA_TEMPR35[17] , \R_DATA_TEMPR36[17] , 
        \R_DATA_TEMPR37[17] , \R_DATA_TEMPR38[17] , 
        \R_DATA_TEMPR39[17] , \R_DATA_TEMPR40[17] , 
        \R_DATA_TEMPR41[17] , \R_DATA_TEMPR42[17] , 
        \R_DATA_TEMPR43[17] , \R_DATA_TEMPR44[17] , 
        \R_DATA_TEMPR45[17] , \R_DATA_TEMPR46[17] , 
        \R_DATA_TEMPR47[17] , \R_DATA_TEMPR48[17] , 
        \R_DATA_TEMPR49[17] , \R_DATA_TEMPR50[17] , 
        \R_DATA_TEMPR51[17] , \R_DATA_TEMPR52[17] , 
        \R_DATA_TEMPR53[17] , \R_DATA_TEMPR54[17] , 
        \R_DATA_TEMPR55[17] , \R_DATA_TEMPR56[17] , 
        \R_DATA_TEMPR57[17] , \R_DATA_TEMPR58[17] , 
        \R_DATA_TEMPR59[17] , \R_DATA_TEMPR60[17] , 
        \R_DATA_TEMPR61[17] , \R_DATA_TEMPR62[17] , 
        \R_DATA_TEMPR63[17] , \R_DATA_TEMPR0[18] , \R_DATA_TEMPR1[18] , 
        \R_DATA_TEMPR2[18] , \R_DATA_TEMPR3[18] , \R_DATA_TEMPR4[18] , 
        \R_DATA_TEMPR5[18] , \R_DATA_TEMPR6[18] , \R_DATA_TEMPR7[18] , 
        \R_DATA_TEMPR8[18] , \R_DATA_TEMPR9[18] , \R_DATA_TEMPR10[18] , 
        \R_DATA_TEMPR11[18] , \R_DATA_TEMPR12[18] , 
        \R_DATA_TEMPR13[18] , \R_DATA_TEMPR14[18] , 
        \R_DATA_TEMPR15[18] , \R_DATA_TEMPR16[18] , 
        \R_DATA_TEMPR17[18] , \R_DATA_TEMPR18[18] , 
        \R_DATA_TEMPR19[18] , \R_DATA_TEMPR20[18] , 
        \R_DATA_TEMPR21[18] , \R_DATA_TEMPR22[18] , 
        \R_DATA_TEMPR23[18] , \R_DATA_TEMPR24[18] , 
        \R_DATA_TEMPR25[18] , \R_DATA_TEMPR26[18] , 
        \R_DATA_TEMPR27[18] , \R_DATA_TEMPR28[18] , 
        \R_DATA_TEMPR29[18] , \R_DATA_TEMPR30[18] , 
        \R_DATA_TEMPR31[18] , \R_DATA_TEMPR32[18] , 
        \R_DATA_TEMPR33[18] , \R_DATA_TEMPR34[18] , 
        \R_DATA_TEMPR35[18] , \R_DATA_TEMPR36[18] , 
        \R_DATA_TEMPR37[18] , \R_DATA_TEMPR38[18] , 
        \R_DATA_TEMPR39[18] , \R_DATA_TEMPR40[18] , 
        \R_DATA_TEMPR41[18] , \R_DATA_TEMPR42[18] , 
        \R_DATA_TEMPR43[18] , \R_DATA_TEMPR44[18] , 
        \R_DATA_TEMPR45[18] , \R_DATA_TEMPR46[18] , 
        \R_DATA_TEMPR47[18] , \R_DATA_TEMPR48[18] , 
        \R_DATA_TEMPR49[18] , \R_DATA_TEMPR50[18] , 
        \R_DATA_TEMPR51[18] , \R_DATA_TEMPR52[18] , 
        \R_DATA_TEMPR53[18] , \R_DATA_TEMPR54[18] , 
        \R_DATA_TEMPR55[18] , \R_DATA_TEMPR56[18] , 
        \R_DATA_TEMPR57[18] , \R_DATA_TEMPR58[18] , 
        \R_DATA_TEMPR59[18] , \R_DATA_TEMPR60[18] , 
        \R_DATA_TEMPR61[18] , \R_DATA_TEMPR62[18] , 
        \R_DATA_TEMPR63[18] , \R_DATA_TEMPR0[19] , \R_DATA_TEMPR1[19] , 
        \R_DATA_TEMPR2[19] , \R_DATA_TEMPR3[19] , \R_DATA_TEMPR4[19] , 
        \R_DATA_TEMPR5[19] , \R_DATA_TEMPR6[19] , \R_DATA_TEMPR7[19] , 
        \R_DATA_TEMPR8[19] , \R_DATA_TEMPR9[19] , \R_DATA_TEMPR10[19] , 
        \R_DATA_TEMPR11[19] , \R_DATA_TEMPR12[19] , 
        \R_DATA_TEMPR13[19] , \R_DATA_TEMPR14[19] , 
        \R_DATA_TEMPR15[19] , \R_DATA_TEMPR16[19] , 
        \R_DATA_TEMPR17[19] , \R_DATA_TEMPR18[19] , 
        \R_DATA_TEMPR19[19] , \R_DATA_TEMPR20[19] , 
        \R_DATA_TEMPR21[19] , \R_DATA_TEMPR22[19] , 
        \R_DATA_TEMPR23[19] , \R_DATA_TEMPR24[19] , 
        \R_DATA_TEMPR25[19] , \R_DATA_TEMPR26[19] , 
        \R_DATA_TEMPR27[19] , \R_DATA_TEMPR28[19] , 
        \R_DATA_TEMPR29[19] , \R_DATA_TEMPR30[19] , 
        \R_DATA_TEMPR31[19] , \R_DATA_TEMPR32[19] , 
        \R_DATA_TEMPR33[19] , \R_DATA_TEMPR34[19] , 
        \R_DATA_TEMPR35[19] , \R_DATA_TEMPR36[19] , 
        \R_DATA_TEMPR37[19] , \R_DATA_TEMPR38[19] , 
        \R_DATA_TEMPR39[19] , \R_DATA_TEMPR40[19] , 
        \R_DATA_TEMPR41[19] , \R_DATA_TEMPR42[19] , 
        \R_DATA_TEMPR43[19] , \R_DATA_TEMPR44[19] , 
        \R_DATA_TEMPR45[19] , \R_DATA_TEMPR46[19] , 
        \R_DATA_TEMPR47[19] , \R_DATA_TEMPR48[19] , 
        \R_DATA_TEMPR49[19] , \R_DATA_TEMPR50[19] , 
        \R_DATA_TEMPR51[19] , \R_DATA_TEMPR52[19] , 
        \R_DATA_TEMPR53[19] , \R_DATA_TEMPR54[19] , 
        \R_DATA_TEMPR55[19] , \R_DATA_TEMPR56[19] , 
        \R_DATA_TEMPR57[19] , \R_DATA_TEMPR58[19] , 
        \R_DATA_TEMPR59[19] , \R_DATA_TEMPR60[19] , 
        \R_DATA_TEMPR61[19] , \R_DATA_TEMPR62[19] , 
        \R_DATA_TEMPR63[19] , \R_DATA_TEMPR0[20] , \R_DATA_TEMPR1[20] , 
        \R_DATA_TEMPR2[20] , \R_DATA_TEMPR3[20] , \R_DATA_TEMPR4[20] , 
        \R_DATA_TEMPR5[20] , \R_DATA_TEMPR6[20] , \R_DATA_TEMPR7[20] , 
        \R_DATA_TEMPR8[20] , \R_DATA_TEMPR9[20] , \R_DATA_TEMPR10[20] , 
        \R_DATA_TEMPR11[20] , \R_DATA_TEMPR12[20] , 
        \R_DATA_TEMPR13[20] , \R_DATA_TEMPR14[20] , 
        \R_DATA_TEMPR15[20] , \R_DATA_TEMPR16[20] , 
        \R_DATA_TEMPR17[20] , \R_DATA_TEMPR18[20] , 
        \R_DATA_TEMPR19[20] , \R_DATA_TEMPR20[20] , 
        \R_DATA_TEMPR21[20] , \R_DATA_TEMPR22[20] , 
        \R_DATA_TEMPR23[20] , \R_DATA_TEMPR24[20] , 
        \R_DATA_TEMPR25[20] , \R_DATA_TEMPR26[20] , 
        \R_DATA_TEMPR27[20] , \R_DATA_TEMPR28[20] , 
        \R_DATA_TEMPR29[20] , \R_DATA_TEMPR30[20] , 
        \R_DATA_TEMPR31[20] , \R_DATA_TEMPR32[20] , 
        \R_DATA_TEMPR33[20] , \R_DATA_TEMPR34[20] , 
        \R_DATA_TEMPR35[20] , \R_DATA_TEMPR36[20] , 
        \R_DATA_TEMPR37[20] , \R_DATA_TEMPR38[20] , 
        \R_DATA_TEMPR39[20] , \R_DATA_TEMPR40[20] , 
        \R_DATA_TEMPR41[20] , \R_DATA_TEMPR42[20] , 
        \R_DATA_TEMPR43[20] , \R_DATA_TEMPR44[20] , 
        \R_DATA_TEMPR45[20] , \R_DATA_TEMPR46[20] , 
        \R_DATA_TEMPR47[20] , \R_DATA_TEMPR48[20] , 
        \R_DATA_TEMPR49[20] , \R_DATA_TEMPR50[20] , 
        \R_DATA_TEMPR51[20] , \R_DATA_TEMPR52[20] , 
        \R_DATA_TEMPR53[20] , \R_DATA_TEMPR54[20] , 
        \R_DATA_TEMPR55[20] , \R_DATA_TEMPR56[20] , 
        \R_DATA_TEMPR57[20] , \R_DATA_TEMPR58[20] , 
        \R_DATA_TEMPR59[20] , \R_DATA_TEMPR60[20] , 
        \R_DATA_TEMPR61[20] , \R_DATA_TEMPR62[20] , 
        \R_DATA_TEMPR63[20] , \R_DATA_TEMPR0[21] , \R_DATA_TEMPR1[21] , 
        \R_DATA_TEMPR2[21] , \R_DATA_TEMPR3[21] , \R_DATA_TEMPR4[21] , 
        \R_DATA_TEMPR5[21] , \R_DATA_TEMPR6[21] , \R_DATA_TEMPR7[21] , 
        \R_DATA_TEMPR8[21] , \R_DATA_TEMPR9[21] , \R_DATA_TEMPR10[21] , 
        \R_DATA_TEMPR11[21] , \R_DATA_TEMPR12[21] , 
        \R_DATA_TEMPR13[21] , \R_DATA_TEMPR14[21] , 
        \R_DATA_TEMPR15[21] , \R_DATA_TEMPR16[21] , 
        \R_DATA_TEMPR17[21] , \R_DATA_TEMPR18[21] , 
        \R_DATA_TEMPR19[21] , \R_DATA_TEMPR20[21] , 
        \R_DATA_TEMPR21[21] , \R_DATA_TEMPR22[21] , 
        \R_DATA_TEMPR23[21] , \R_DATA_TEMPR24[21] , 
        \R_DATA_TEMPR25[21] , \R_DATA_TEMPR26[21] , 
        \R_DATA_TEMPR27[21] , \R_DATA_TEMPR28[21] , 
        \R_DATA_TEMPR29[21] , \R_DATA_TEMPR30[21] , 
        \R_DATA_TEMPR31[21] , \R_DATA_TEMPR32[21] , 
        \R_DATA_TEMPR33[21] , \R_DATA_TEMPR34[21] , 
        \R_DATA_TEMPR35[21] , \R_DATA_TEMPR36[21] , 
        \R_DATA_TEMPR37[21] , \R_DATA_TEMPR38[21] , 
        \R_DATA_TEMPR39[21] , \R_DATA_TEMPR40[21] , 
        \R_DATA_TEMPR41[21] , \R_DATA_TEMPR42[21] , 
        \R_DATA_TEMPR43[21] , \R_DATA_TEMPR44[21] , 
        \R_DATA_TEMPR45[21] , \R_DATA_TEMPR46[21] , 
        \R_DATA_TEMPR47[21] , \R_DATA_TEMPR48[21] , 
        \R_DATA_TEMPR49[21] , \R_DATA_TEMPR50[21] , 
        \R_DATA_TEMPR51[21] , \R_DATA_TEMPR52[21] , 
        \R_DATA_TEMPR53[21] , \R_DATA_TEMPR54[21] , 
        \R_DATA_TEMPR55[21] , \R_DATA_TEMPR56[21] , 
        \R_DATA_TEMPR57[21] , \R_DATA_TEMPR58[21] , 
        \R_DATA_TEMPR59[21] , \R_DATA_TEMPR60[21] , 
        \R_DATA_TEMPR61[21] , \R_DATA_TEMPR62[21] , 
        \R_DATA_TEMPR63[21] , \R_DATA_TEMPR0[22] , \R_DATA_TEMPR1[22] , 
        \R_DATA_TEMPR2[22] , \R_DATA_TEMPR3[22] , \R_DATA_TEMPR4[22] , 
        \R_DATA_TEMPR5[22] , \R_DATA_TEMPR6[22] , \R_DATA_TEMPR7[22] , 
        \R_DATA_TEMPR8[22] , \R_DATA_TEMPR9[22] , \R_DATA_TEMPR10[22] , 
        \R_DATA_TEMPR11[22] , \R_DATA_TEMPR12[22] , 
        \R_DATA_TEMPR13[22] , \R_DATA_TEMPR14[22] , 
        \R_DATA_TEMPR15[22] , \R_DATA_TEMPR16[22] , 
        \R_DATA_TEMPR17[22] , \R_DATA_TEMPR18[22] , 
        \R_DATA_TEMPR19[22] , \R_DATA_TEMPR20[22] , 
        \R_DATA_TEMPR21[22] , \R_DATA_TEMPR22[22] , 
        \R_DATA_TEMPR23[22] , \R_DATA_TEMPR24[22] , 
        \R_DATA_TEMPR25[22] , \R_DATA_TEMPR26[22] , 
        \R_DATA_TEMPR27[22] , \R_DATA_TEMPR28[22] , 
        \R_DATA_TEMPR29[22] , \R_DATA_TEMPR30[22] , 
        \R_DATA_TEMPR31[22] , \R_DATA_TEMPR32[22] , 
        \R_DATA_TEMPR33[22] , \R_DATA_TEMPR34[22] , 
        \R_DATA_TEMPR35[22] , \R_DATA_TEMPR36[22] , 
        \R_DATA_TEMPR37[22] , \R_DATA_TEMPR38[22] , 
        \R_DATA_TEMPR39[22] , \R_DATA_TEMPR40[22] , 
        \R_DATA_TEMPR41[22] , \R_DATA_TEMPR42[22] , 
        \R_DATA_TEMPR43[22] , \R_DATA_TEMPR44[22] , 
        \R_DATA_TEMPR45[22] , \R_DATA_TEMPR46[22] , 
        \R_DATA_TEMPR47[22] , \R_DATA_TEMPR48[22] , 
        \R_DATA_TEMPR49[22] , \R_DATA_TEMPR50[22] , 
        \R_DATA_TEMPR51[22] , \R_DATA_TEMPR52[22] , 
        \R_DATA_TEMPR53[22] , \R_DATA_TEMPR54[22] , 
        \R_DATA_TEMPR55[22] , \R_DATA_TEMPR56[22] , 
        \R_DATA_TEMPR57[22] , \R_DATA_TEMPR58[22] , 
        \R_DATA_TEMPR59[22] , \R_DATA_TEMPR60[22] , 
        \R_DATA_TEMPR61[22] , \R_DATA_TEMPR62[22] , 
        \R_DATA_TEMPR63[22] , \R_DATA_TEMPR0[23] , \R_DATA_TEMPR1[23] , 
        \R_DATA_TEMPR2[23] , \R_DATA_TEMPR3[23] , \R_DATA_TEMPR4[23] , 
        \R_DATA_TEMPR5[23] , \R_DATA_TEMPR6[23] , \R_DATA_TEMPR7[23] , 
        \R_DATA_TEMPR8[23] , \R_DATA_TEMPR9[23] , \R_DATA_TEMPR10[23] , 
        \R_DATA_TEMPR11[23] , \R_DATA_TEMPR12[23] , 
        \R_DATA_TEMPR13[23] , \R_DATA_TEMPR14[23] , 
        \R_DATA_TEMPR15[23] , \R_DATA_TEMPR16[23] , 
        \R_DATA_TEMPR17[23] , \R_DATA_TEMPR18[23] , 
        \R_DATA_TEMPR19[23] , \R_DATA_TEMPR20[23] , 
        \R_DATA_TEMPR21[23] , \R_DATA_TEMPR22[23] , 
        \R_DATA_TEMPR23[23] , \R_DATA_TEMPR24[23] , 
        \R_DATA_TEMPR25[23] , \R_DATA_TEMPR26[23] , 
        \R_DATA_TEMPR27[23] , \R_DATA_TEMPR28[23] , 
        \R_DATA_TEMPR29[23] , \R_DATA_TEMPR30[23] , 
        \R_DATA_TEMPR31[23] , \R_DATA_TEMPR32[23] , 
        \R_DATA_TEMPR33[23] , \R_DATA_TEMPR34[23] , 
        \R_DATA_TEMPR35[23] , \R_DATA_TEMPR36[23] , 
        \R_DATA_TEMPR37[23] , \R_DATA_TEMPR38[23] , 
        \R_DATA_TEMPR39[23] , \R_DATA_TEMPR40[23] , 
        \R_DATA_TEMPR41[23] , \R_DATA_TEMPR42[23] , 
        \R_DATA_TEMPR43[23] , \R_DATA_TEMPR44[23] , 
        \R_DATA_TEMPR45[23] , \R_DATA_TEMPR46[23] , 
        \R_DATA_TEMPR47[23] , \R_DATA_TEMPR48[23] , 
        \R_DATA_TEMPR49[23] , \R_DATA_TEMPR50[23] , 
        \R_DATA_TEMPR51[23] , \R_DATA_TEMPR52[23] , 
        \R_DATA_TEMPR53[23] , \R_DATA_TEMPR54[23] , 
        \R_DATA_TEMPR55[23] , \R_DATA_TEMPR56[23] , 
        \R_DATA_TEMPR57[23] , \R_DATA_TEMPR58[23] , 
        \R_DATA_TEMPR59[23] , \R_DATA_TEMPR60[23] , 
        \R_DATA_TEMPR61[23] , \R_DATA_TEMPR62[23] , 
        \R_DATA_TEMPR63[23] , \R_DATA_TEMPR0[24] , \R_DATA_TEMPR1[24] , 
        \R_DATA_TEMPR2[24] , \R_DATA_TEMPR3[24] , \R_DATA_TEMPR4[24] , 
        \R_DATA_TEMPR5[24] , \R_DATA_TEMPR6[24] , \R_DATA_TEMPR7[24] , 
        \R_DATA_TEMPR8[24] , \R_DATA_TEMPR9[24] , \R_DATA_TEMPR10[24] , 
        \R_DATA_TEMPR11[24] , \R_DATA_TEMPR12[24] , 
        \R_DATA_TEMPR13[24] , \R_DATA_TEMPR14[24] , 
        \R_DATA_TEMPR15[24] , \R_DATA_TEMPR16[24] , 
        \R_DATA_TEMPR17[24] , \R_DATA_TEMPR18[24] , 
        \R_DATA_TEMPR19[24] , \R_DATA_TEMPR20[24] , 
        \R_DATA_TEMPR21[24] , \R_DATA_TEMPR22[24] , 
        \R_DATA_TEMPR23[24] , \R_DATA_TEMPR24[24] , 
        \R_DATA_TEMPR25[24] , \R_DATA_TEMPR26[24] , 
        \R_DATA_TEMPR27[24] , \R_DATA_TEMPR28[24] , 
        \R_DATA_TEMPR29[24] , \R_DATA_TEMPR30[24] , 
        \R_DATA_TEMPR31[24] , \R_DATA_TEMPR32[24] , 
        \R_DATA_TEMPR33[24] , \R_DATA_TEMPR34[24] , 
        \R_DATA_TEMPR35[24] , \R_DATA_TEMPR36[24] , 
        \R_DATA_TEMPR37[24] , \R_DATA_TEMPR38[24] , 
        \R_DATA_TEMPR39[24] , \R_DATA_TEMPR40[24] , 
        \R_DATA_TEMPR41[24] , \R_DATA_TEMPR42[24] , 
        \R_DATA_TEMPR43[24] , \R_DATA_TEMPR44[24] , 
        \R_DATA_TEMPR45[24] , \R_DATA_TEMPR46[24] , 
        \R_DATA_TEMPR47[24] , \R_DATA_TEMPR48[24] , 
        \R_DATA_TEMPR49[24] , \R_DATA_TEMPR50[24] , 
        \R_DATA_TEMPR51[24] , \R_DATA_TEMPR52[24] , 
        \R_DATA_TEMPR53[24] , \R_DATA_TEMPR54[24] , 
        \R_DATA_TEMPR55[24] , \R_DATA_TEMPR56[24] , 
        \R_DATA_TEMPR57[24] , \R_DATA_TEMPR58[24] , 
        \R_DATA_TEMPR59[24] , \R_DATA_TEMPR60[24] , 
        \R_DATA_TEMPR61[24] , \R_DATA_TEMPR62[24] , 
        \R_DATA_TEMPR63[24] , \R_DATA_TEMPR0[25] , \R_DATA_TEMPR1[25] , 
        \R_DATA_TEMPR2[25] , \R_DATA_TEMPR3[25] , \R_DATA_TEMPR4[25] , 
        \R_DATA_TEMPR5[25] , \R_DATA_TEMPR6[25] , \R_DATA_TEMPR7[25] , 
        \R_DATA_TEMPR8[25] , \R_DATA_TEMPR9[25] , \R_DATA_TEMPR10[25] , 
        \R_DATA_TEMPR11[25] , \R_DATA_TEMPR12[25] , 
        \R_DATA_TEMPR13[25] , \R_DATA_TEMPR14[25] , 
        \R_DATA_TEMPR15[25] , \R_DATA_TEMPR16[25] , 
        \R_DATA_TEMPR17[25] , \R_DATA_TEMPR18[25] , 
        \R_DATA_TEMPR19[25] , \R_DATA_TEMPR20[25] , 
        \R_DATA_TEMPR21[25] , \R_DATA_TEMPR22[25] , 
        \R_DATA_TEMPR23[25] , \R_DATA_TEMPR24[25] , 
        \R_DATA_TEMPR25[25] , \R_DATA_TEMPR26[25] , 
        \R_DATA_TEMPR27[25] , \R_DATA_TEMPR28[25] , 
        \R_DATA_TEMPR29[25] , \R_DATA_TEMPR30[25] , 
        \R_DATA_TEMPR31[25] , \R_DATA_TEMPR32[25] , 
        \R_DATA_TEMPR33[25] , \R_DATA_TEMPR34[25] , 
        \R_DATA_TEMPR35[25] , \R_DATA_TEMPR36[25] , 
        \R_DATA_TEMPR37[25] , \R_DATA_TEMPR38[25] , 
        \R_DATA_TEMPR39[25] , \R_DATA_TEMPR40[25] , 
        \R_DATA_TEMPR41[25] , \R_DATA_TEMPR42[25] , 
        \R_DATA_TEMPR43[25] , \R_DATA_TEMPR44[25] , 
        \R_DATA_TEMPR45[25] , \R_DATA_TEMPR46[25] , 
        \R_DATA_TEMPR47[25] , \R_DATA_TEMPR48[25] , 
        \R_DATA_TEMPR49[25] , \R_DATA_TEMPR50[25] , 
        \R_DATA_TEMPR51[25] , \R_DATA_TEMPR52[25] , 
        \R_DATA_TEMPR53[25] , \R_DATA_TEMPR54[25] , 
        \R_DATA_TEMPR55[25] , \R_DATA_TEMPR56[25] , 
        \R_DATA_TEMPR57[25] , \R_DATA_TEMPR58[25] , 
        \R_DATA_TEMPR59[25] , \R_DATA_TEMPR60[25] , 
        \R_DATA_TEMPR61[25] , \R_DATA_TEMPR62[25] , 
        \R_DATA_TEMPR63[25] , \R_DATA_TEMPR0[26] , \R_DATA_TEMPR1[26] , 
        \R_DATA_TEMPR2[26] , \R_DATA_TEMPR3[26] , \R_DATA_TEMPR4[26] , 
        \R_DATA_TEMPR5[26] , \R_DATA_TEMPR6[26] , \R_DATA_TEMPR7[26] , 
        \R_DATA_TEMPR8[26] , \R_DATA_TEMPR9[26] , \R_DATA_TEMPR10[26] , 
        \R_DATA_TEMPR11[26] , \R_DATA_TEMPR12[26] , 
        \R_DATA_TEMPR13[26] , \R_DATA_TEMPR14[26] , 
        \R_DATA_TEMPR15[26] , \R_DATA_TEMPR16[26] , 
        \R_DATA_TEMPR17[26] , \R_DATA_TEMPR18[26] , 
        \R_DATA_TEMPR19[26] , \R_DATA_TEMPR20[26] , 
        \R_DATA_TEMPR21[26] , \R_DATA_TEMPR22[26] , 
        \R_DATA_TEMPR23[26] , \R_DATA_TEMPR24[26] , 
        \R_DATA_TEMPR25[26] , \R_DATA_TEMPR26[26] , 
        \R_DATA_TEMPR27[26] , \R_DATA_TEMPR28[26] , 
        \R_DATA_TEMPR29[26] , \R_DATA_TEMPR30[26] , 
        \R_DATA_TEMPR31[26] , \R_DATA_TEMPR32[26] , 
        \R_DATA_TEMPR33[26] , \R_DATA_TEMPR34[26] , 
        \R_DATA_TEMPR35[26] , \R_DATA_TEMPR36[26] , 
        \R_DATA_TEMPR37[26] , \R_DATA_TEMPR38[26] , 
        \R_DATA_TEMPR39[26] , \R_DATA_TEMPR40[26] , 
        \R_DATA_TEMPR41[26] , \R_DATA_TEMPR42[26] , 
        \R_DATA_TEMPR43[26] , \R_DATA_TEMPR44[26] , 
        \R_DATA_TEMPR45[26] , \R_DATA_TEMPR46[26] , 
        \R_DATA_TEMPR47[26] , \R_DATA_TEMPR48[26] , 
        \R_DATA_TEMPR49[26] , \R_DATA_TEMPR50[26] , 
        \R_DATA_TEMPR51[26] , \R_DATA_TEMPR52[26] , 
        \R_DATA_TEMPR53[26] , \R_DATA_TEMPR54[26] , 
        \R_DATA_TEMPR55[26] , \R_DATA_TEMPR56[26] , 
        \R_DATA_TEMPR57[26] , \R_DATA_TEMPR58[26] , 
        \R_DATA_TEMPR59[26] , \R_DATA_TEMPR60[26] , 
        \R_DATA_TEMPR61[26] , \R_DATA_TEMPR62[26] , 
        \R_DATA_TEMPR63[26] , \R_DATA_TEMPR0[27] , \R_DATA_TEMPR1[27] , 
        \R_DATA_TEMPR2[27] , \R_DATA_TEMPR3[27] , \R_DATA_TEMPR4[27] , 
        \R_DATA_TEMPR5[27] , \R_DATA_TEMPR6[27] , \R_DATA_TEMPR7[27] , 
        \R_DATA_TEMPR8[27] , \R_DATA_TEMPR9[27] , \R_DATA_TEMPR10[27] , 
        \R_DATA_TEMPR11[27] , \R_DATA_TEMPR12[27] , 
        \R_DATA_TEMPR13[27] , \R_DATA_TEMPR14[27] , 
        \R_DATA_TEMPR15[27] , \R_DATA_TEMPR16[27] , 
        \R_DATA_TEMPR17[27] , \R_DATA_TEMPR18[27] , 
        \R_DATA_TEMPR19[27] , \R_DATA_TEMPR20[27] , 
        \R_DATA_TEMPR21[27] , \R_DATA_TEMPR22[27] , 
        \R_DATA_TEMPR23[27] , \R_DATA_TEMPR24[27] , 
        \R_DATA_TEMPR25[27] , \R_DATA_TEMPR26[27] , 
        \R_DATA_TEMPR27[27] , \R_DATA_TEMPR28[27] , 
        \R_DATA_TEMPR29[27] , \R_DATA_TEMPR30[27] , 
        \R_DATA_TEMPR31[27] , \R_DATA_TEMPR32[27] , 
        \R_DATA_TEMPR33[27] , \R_DATA_TEMPR34[27] , 
        \R_DATA_TEMPR35[27] , \R_DATA_TEMPR36[27] , 
        \R_DATA_TEMPR37[27] , \R_DATA_TEMPR38[27] , 
        \R_DATA_TEMPR39[27] , \R_DATA_TEMPR40[27] , 
        \R_DATA_TEMPR41[27] , \R_DATA_TEMPR42[27] , 
        \R_DATA_TEMPR43[27] , \R_DATA_TEMPR44[27] , 
        \R_DATA_TEMPR45[27] , \R_DATA_TEMPR46[27] , 
        \R_DATA_TEMPR47[27] , \R_DATA_TEMPR48[27] , 
        \R_DATA_TEMPR49[27] , \R_DATA_TEMPR50[27] , 
        \R_DATA_TEMPR51[27] , \R_DATA_TEMPR52[27] , 
        \R_DATA_TEMPR53[27] , \R_DATA_TEMPR54[27] , 
        \R_DATA_TEMPR55[27] , \R_DATA_TEMPR56[27] , 
        \R_DATA_TEMPR57[27] , \R_DATA_TEMPR58[27] , 
        \R_DATA_TEMPR59[27] , \R_DATA_TEMPR60[27] , 
        \R_DATA_TEMPR61[27] , \R_DATA_TEMPR62[27] , 
        \R_DATA_TEMPR63[27] , \R_DATA_TEMPR0[28] , \R_DATA_TEMPR1[28] , 
        \R_DATA_TEMPR2[28] , \R_DATA_TEMPR3[28] , \R_DATA_TEMPR4[28] , 
        \R_DATA_TEMPR5[28] , \R_DATA_TEMPR6[28] , \R_DATA_TEMPR7[28] , 
        \R_DATA_TEMPR8[28] , \R_DATA_TEMPR9[28] , \R_DATA_TEMPR10[28] , 
        \R_DATA_TEMPR11[28] , \R_DATA_TEMPR12[28] , 
        \R_DATA_TEMPR13[28] , \R_DATA_TEMPR14[28] , 
        \R_DATA_TEMPR15[28] , \R_DATA_TEMPR16[28] , 
        \R_DATA_TEMPR17[28] , \R_DATA_TEMPR18[28] , 
        \R_DATA_TEMPR19[28] , \R_DATA_TEMPR20[28] , 
        \R_DATA_TEMPR21[28] , \R_DATA_TEMPR22[28] , 
        \R_DATA_TEMPR23[28] , \R_DATA_TEMPR24[28] , 
        \R_DATA_TEMPR25[28] , \R_DATA_TEMPR26[28] , 
        \R_DATA_TEMPR27[28] , \R_DATA_TEMPR28[28] , 
        \R_DATA_TEMPR29[28] , \R_DATA_TEMPR30[28] , 
        \R_DATA_TEMPR31[28] , \R_DATA_TEMPR32[28] , 
        \R_DATA_TEMPR33[28] , \R_DATA_TEMPR34[28] , 
        \R_DATA_TEMPR35[28] , \R_DATA_TEMPR36[28] , 
        \R_DATA_TEMPR37[28] , \R_DATA_TEMPR38[28] , 
        \R_DATA_TEMPR39[28] , \R_DATA_TEMPR40[28] , 
        \R_DATA_TEMPR41[28] , \R_DATA_TEMPR42[28] , 
        \R_DATA_TEMPR43[28] , \R_DATA_TEMPR44[28] , 
        \R_DATA_TEMPR45[28] , \R_DATA_TEMPR46[28] , 
        \R_DATA_TEMPR47[28] , \R_DATA_TEMPR48[28] , 
        \R_DATA_TEMPR49[28] , \R_DATA_TEMPR50[28] , 
        \R_DATA_TEMPR51[28] , \R_DATA_TEMPR52[28] , 
        \R_DATA_TEMPR53[28] , \R_DATA_TEMPR54[28] , 
        \R_DATA_TEMPR55[28] , \R_DATA_TEMPR56[28] , 
        \R_DATA_TEMPR57[28] , \R_DATA_TEMPR58[28] , 
        \R_DATA_TEMPR59[28] , \R_DATA_TEMPR60[28] , 
        \R_DATA_TEMPR61[28] , \R_DATA_TEMPR62[28] , 
        \R_DATA_TEMPR63[28] , \R_DATA_TEMPR0[29] , \R_DATA_TEMPR1[29] , 
        \R_DATA_TEMPR2[29] , \R_DATA_TEMPR3[29] , \R_DATA_TEMPR4[29] , 
        \R_DATA_TEMPR5[29] , \R_DATA_TEMPR6[29] , \R_DATA_TEMPR7[29] , 
        \R_DATA_TEMPR8[29] , \R_DATA_TEMPR9[29] , \R_DATA_TEMPR10[29] , 
        \R_DATA_TEMPR11[29] , \R_DATA_TEMPR12[29] , 
        \R_DATA_TEMPR13[29] , \R_DATA_TEMPR14[29] , 
        \R_DATA_TEMPR15[29] , \R_DATA_TEMPR16[29] , 
        \R_DATA_TEMPR17[29] , \R_DATA_TEMPR18[29] , 
        \R_DATA_TEMPR19[29] , \R_DATA_TEMPR20[29] , 
        \R_DATA_TEMPR21[29] , \R_DATA_TEMPR22[29] , 
        \R_DATA_TEMPR23[29] , \R_DATA_TEMPR24[29] , 
        \R_DATA_TEMPR25[29] , \R_DATA_TEMPR26[29] , 
        \R_DATA_TEMPR27[29] , \R_DATA_TEMPR28[29] , 
        \R_DATA_TEMPR29[29] , \R_DATA_TEMPR30[29] , 
        \R_DATA_TEMPR31[29] , \R_DATA_TEMPR32[29] , 
        \R_DATA_TEMPR33[29] , \R_DATA_TEMPR34[29] , 
        \R_DATA_TEMPR35[29] , \R_DATA_TEMPR36[29] , 
        \R_DATA_TEMPR37[29] , \R_DATA_TEMPR38[29] , 
        \R_DATA_TEMPR39[29] , \R_DATA_TEMPR40[29] , 
        \R_DATA_TEMPR41[29] , \R_DATA_TEMPR42[29] , 
        \R_DATA_TEMPR43[29] , \R_DATA_TEMPR44[29] , 
        \R_DATA_TEMPR45[29] , \R_DATA_TEMPR46[29] , 
        \R_DATA_TEMPR47[29] , \R_DATA_TEMPR48[29] , 
        \R_DATA_TEMPR49[29] , \R_DATA_TEMPR50[29] , 
        \R_DATA_TEMPR51[29] , \R_DATA_TEMPR52[29] , 
        \R_DATA_TEMPR53[29] , \R_DATA_TEMPR54[29] , 
        \R_DATA_TEMPR55[29] , \R_DATA_TEMPR56[29] , 
        \R_DATA_TEMPR57[29] , \R_DATA_TEMPR58[29] , 
        \R_DATA_TEMPR59[29] , \R_DATA_TEMPR60[29] , 
        \R_DATA_TEMPR61[29] , \R_DATA_TEMPR62[29] , 
        \R_DATA_TEMPR63[29] , \R_DATA_TEMPR0[30] , \R_DATA_TEMPR1[30] , 
        \R_DATA_TEMPR2[30] , \R_DATA_TEMPR3[30] , \R_DATA_TEMPR4[30] , 
        \R_DATA_TEMPR5[30] , \R_DATA_TEMPR6[30] , \R_DATA_TEMPR7[30] , 
        \R_DATA_TEMPR8[30] , \R_DATA_TEMPR9[30] , \R_DATA_TEMPR10[30] , 
        \R_DATA_TEMPR11[30] , \R_DATA_TEMPR12[30] , 
        \R_DATA_TEMPR13[30] , \R_DATA_TEMPR14[30] , 
        \R_DATA_TEMPR15[30] , \R_DATA_TEMPR16[30] , 
        \R_DATA_TEMPR17[30] , \R_DATA_TEMPR18[30] , 
        \R_DATA_TEMPR19[30] , \R_DATA_TEMPR20[30] , 
        \R_DATA_TEMPR21[30] , \R_DATA_TEMPR22[30] , 
        \R_DATA_TEMPR23[30] , \R_DATA_TEMPR24[30] , 
        \R_DATA_TEMPR25[30] , \R_DATA_TEMPR26[30] , 
        \R_DATA_TEMPR27[30] , \R_DATA_TEMPR28[30] , 
        \R_DATA_TEMPR29[30] , \R_DATA_TEMPR30[30] , 
        \R_DATA_TEMPR31[30] , \R_DATA_TEMPR32[30] , 
        \R_DATA_TEMPR33[30] , \R_DATA_TEMPR34[30] , 
        \R_DATA_TEMPR35[30] , \R_DATA_TEMPR36[30] , 
        \R_DATA_TEMPR37[30] , \R_DATA_TEMPR38[30] , 
        \R_DATA_TEMPR39[30] , \R_DATA_TEMPR40[30] , 
        \R_DATA_TEMPR41[30] , \R_DATA_TEMPR42[30] , 
        \R_DATA_TEMPR43[30] , \R_DATA_TEMPR44[30] , 
        \R_DATA_TEMPR45[30] , \R_DATA_TEMPR46[30] , 
        \R_DATA_TEMPR47[30] , \R_DATA_TEMPR48[30] , 
        \R_DATA_TEMPR49[30] , \R_DATA_TEMPR50[30] , 
        \R_DATA_TEMPR51[30] , \R_DATA_TEMPR52[30] , 
        \R_DATA_TEMPR53[30] , \R_DATA_TEMPR54[30] , 
        \R_DATA_TEMPR55[30] , \R_DATA_TEMPR56[30] , 
        \R_DATA_TEMPR57[30] , \R_DATA_TEMPR58[30] , 
        \R_DATA_TEMPR59[30] , \R_DATA_TEMPR60[30] , 
        \R_DATA_TEMPR61[30] , \R_DATA_TEMPR62[30] , 
        \R_DATA_TEMPR63[30] , \R_DATA_TEMPR0[31] , \R_DATA_TEMPR1[31] , 
        \R_DATA_TEMPR2[31] , \R_DATA_TEMPR3[31] , \R_DATA_TEMPR4[31] , 
        \R_DATA_TEMPR5[31] , \R_DATA_TEMPR6[31] , \R_DATA_TEMPR7[31] , 
        \R_DATA_TEMPR8[31] , \R_DATA_TEMPR9[31] , \R_DATA_TEMPR10[31] , 
        \R_DATA_TEMPR11[31] , \R_DATA_TEMPR12[31] , 
        \R_DATA_TEMPR13[31] , \R_DATA_TEMPR14[31] , 
        \R_DATA_TEMPR15[31] , \R_DATA_TEMPR16[31] , 
        \R_DATA_TEMPR17[31] , \R_DATA_TEMPR18[31] , 
        \R_DATA_TEMPR19[31] , \R_DATA_TEMPR20[31] , 
        \R_DATA_TEMPR21[31] , \R_DATA_TEMPR22[31] , 
        \R_DATA_TEMPR23[31] , \R_DATA_TEMPR24[31] , 
        \R_DATA_TEMPR25[31] , \R_DATA_TEMPR26[31] , 
        \R_DATA_TEMPR27[31] , \R_DATA_TEMPR28[31] , 
        \R_DATA_TEMPR29[31] , \R_DATA_TEMPR30[31] , 
        \R_DATA_TEMPR31[31] , \R_DATA_TEMPR32[31] , 
        \R_DATA_TEMPR33[31] , \R_DATA_TEMPR34[31] , 
        \R_DATA_TEMPR35[31] , \R_DATA_TEMPR36[31] , 
        \R_DATA_TEMPR37[31] , \R_DATA_TEMPR38[31] , 
        \R_DATA_TEMPR39[31] , \R_DATA_TEMPR40[31] , 
        \R_DATA_TEMPR41[31] , \R_DATA_TEMPR42[31] , 
        \R_DATA_TEMPR43[31] , \R_DATA_TEMPR44[31] , 
        \R_DATA_TEMPR45[31] , \R_DATA_TEMPR46[31] , 
        \R_DATA_TEMPR47[31] , \R_DATA_TEMPR48[31] , 
        \R_DATA_TEMPR49[31] , \R_DATA_TEMPR50[31] , 
        \R_DATA_TEMPR51[31] , \R_DATA_TEMPR52[31] , 
        \R_DATA_TEMPR53[31] , \R_DATA_TEMPR54[31] , 
        \R_DATA_TEMPR55[31] , \R_DATA_TEMPR56[31] , 
        \R_DATA_TEMPR57[31] , \R_DATA_TEMPR58[31] , 
        \R_DATA_TEMPR59[31] , \R_DATA_TEMPR60[31] , 
        \R_DATA_TEMPR61[31] , \R_DATA_TEMPR62[31] , 
        \R_DATA_TEMPR63[31] , \R_DATA_TEMPR0[32] , \R_DATA_TEMPR1[32] , 
        \R_DATA_TEMPR2[32] , \R_DATA_TEMPR3[32] , \R_DATA_TEMPR4[32] , 
        \R_DATA_TEMPR5[32] , \R_DATA_TEMPR6[32] , \R_DATA_TEMPR7[32] , 
        \R_DATA_TEMPR8[32] , \R_DATA_TEMPR9[32] , \R_DATA_TEMPR10[32] , 
        \R_DATA_TEMPR11[32] , \R_DATA_TEMPR12[32] , 
        \R_DATA_TEMPR13[32] , \R_DATA_TEMPR14[32] , 
        \R_DATA_TEMPR15[32] , \R_DATA_TEMPR16[32] , 
        \R_DATA_TEMPR17[32] , \R_DATA_TEMPR18[32] , 
        \R_DATA_TEMPR19[32] , \R_DATA_TEMPR20[32] , 
        \R_DATA_TEMPR21[32] , \R_DATA_TEMPR22[32] , 
        \R_DATA_TEMPR23[32] , \R_DATA_TEMPR24[32] , 
        \R_DATA_TEMPR25[32] , \R_DATA_TEMPR26[32] , 
        \R_DATA_TEMPR27[32] , \R_DATA_TEMPR28[32] , 
        \R_DATA_TEMPR29[32] , \R_DATA_TEMPR30[32] , 
        \R_DATA_TEMPR31[32] , \R_DATA_TEMPR32[32] , 
        \R_DATA_TEMPR33[32] , \R_DATA_TEMPR34[32] , 
        \R_DATA_TEMPR35[32] , \R_DATA_TEMPR36[32] , 
        \R_DATA_TEMPR37[32] , \R_DATA_TEMPR38[32] , 
        \R_DATA_TEMPR39[32] , \R_DATA_TEMPR40[32] , 
        \R_DATA_TEMPR41[32] , \R_DATA_TEMPR42[32] , 
        \R_DATA_TEMPR43[32] , \R_DATA_TEMPR44[32] , 
        \R_DATA_TEMPR45[32] , \R_DATA_TEMPR46[32] , 
        \R_DATA_TEMPR47[32] , \R_DATA_TEMPR48[32] , 
        \R_DATA_TEMPR49[32] , \R_DATA_TEMPR50[32] , 
        \R_DATA_TEMPR51[32] , \R_DATA_TEMPR52[32] , 
        \R_DATA_TEMPR53[32] , \R_DATA_TEMPR54[32] , 
        \R_DATA_TEMPR55[32] , \R_DATA_TEMPR56[32] , 
        \R_DATA_TEMPR57[32] , \R_DATA_TEMPR58[32] , 
        \R_DATA_TEMPR59[32] , \R_DATA_TEMPR60[32] , 
        \R_DATA_TEMPR61[32] , \R_DATA_TEMPR62[32] , 
        \R_DATA_TEMPR63[32] , \R_DATA_TEMPR0[33] , \R_DATA_TEMPR1[33] , 
        \R_DATA_TEMPR2[33] , \R_DATA_TEMPR3[33] , \R_DATA_TEMPR4[33] , 
        \R_DATA_TEMPR5[33] , \R_DATA_TEMPR6[33] , \R_DATA_TEMPR7[33] , 
        \R_DATA_TEMPR8[33] , \R_DATA_TEMPR9[33] , \R_DATA_TEMPR10[33] , 
        \R_DATA_TEMPR11[33] , \R_DATA_TEMPR12[33] , 
        \R_DATA_TEMPR13[33] , \R_DATA_TEMPR14[33] , 
        \R_DATA_TEMPR15[33] , \R_DATA_TEMPR16[33] , 
        \R_DATA_TEMPR17[33] , \R_DATA_TEMPR18[33] , 
        \R_DATA_TEMPR19[33] , \R_DATA_TEMPR20[33] , 
        \R_DATA_TEMPR21[33] , \R_DATA_TEMPR22[33] , 
        \R_DATA_TEMPR23[33] , \R_DATA_TEMPR24[33] , 
        \R_DATA_TEMPR25[33] , \R_DATA_TEMPR26[33] , 
        \R_DATA_TEMPR27[33] , \R_DATA_TEMPR28[33] , 
        \R_DATA_TEMPR29[33] , \R_DATA_TEMPR30[33] , 
        \R_DATA_TEMPR31[33] , \R_DATA_TEMPR32[33] , 
        \R_DATA_TEMPR33[33] , \R_DATA_TEMPR34[33] , 
        \R_DATA_TEMPR35[33] , \R_DATA_TEMPR36[33] , 
        \R_DATA_TEMPR37[33] , \R_DATA_TEMPR38[33] , 
        \R_DATA_TEMPR39[33] , \R_DATA_TEMPR40[33] , 
        \R_DATA_TEMPR41[33] , \R_DATA_TEMPR42[33] , 
        \R_DATA_TEMPR43[33] , \R_DATA_TEMPR44[33] , 
        \R_DATA_TEMPR45[33] , \R_DATA_TEMPR46[33] , 
        \R_DATA_TEMPR47[33] , \R_DATA_TEMPR48[33] , 
        \R_DATA_TEMPR49[33] , \R_DATA_TEMPR50[33] , 
        \R_DATA_TEMPR51[33] , \R_DATA_TEMPR52[33] , 
        \R_DATA_TEMPR53[33] , \R_DATA_TEMPR54[33] , 
        \R_DATA_TEMPR55[33] , \R_DATA_TEMPR56[33] , 
        \R_DATA_TEMPR57[33] , \R_DATA_TEMPR58[33] , 
        \R_DATA_TEMPR59[33] , \R_DATA_TEMPR60[33] , 
        \R_DATA_TEMPR61[33] , \R_DATA_TEMPR62[33] , 
        \R_DATA_TEMPR63[33] , \R_DATA_TEMPR0[34] , \R_DATA_TEMPR1[34] , 
        \R_DATA_TEMPR2[34] , \R_DATA_TEMPR3[34] , \R_DATA_TEMPR4[34] , 
        \R_DATA_TEMPR5[34] , \R_DATA_TEMPR6[34] , \R_DATA_TEMPR7[34] , 
        \R_DATA_TEMPR8[34] , \R_DATA_TEMPR9[34] , \R_DATA_TEMPR10[34] , 
        \R_DATA_TEMPR11[34] , \R_DATA_TEMPR12[34] , 
        \R_DATA_TEMPR13[34] , \R_DATA_TEMPR14[34] , 
        \R_DATA_TEMPR15[34] , \R_DATA_TEMPR16[34] , 
        \R_DATA_TEMPR17[34] , \R_DATA_TEMPR18[34] , 
        \R_DATA_TEMPR19[34] , \R_DATA_TEMPR20[34] , 
        \R_DATA_TEMPR21[34] , \R_DATA_TEMPR22[34] , 
        \R_DATA_TEMPR23[34] , \R_DATA_TEMPR24[34] , 
        \R_DATA_TEMPR25[34] , \R_DATA_TEMPR26[34] , 
        \R_DATA_TEMPR27[34] , \R_DATA_TEMPR28[34] , 
        \R_DATA_TEMPR29[34] , \R_DATA_TEMPR30[34] , 
        \R_DATA_TEMPR31[34] , \R_DATA_TEMPR32[34] , 
        \R_DATA_TEMPR33[34] , \R_DATA_TEMPR34[34] , 
        \R_DATA_TEMPR35[34] , \R_DATA_TEMPR36[34] , 
        \R_DATA_TEMPR37[34] , \R_DATA_TEMPR38[34] , 
        \R_DATA_TEMPR39[34] , \R_DATA_TEMPR40[34] , 
        \R_DATA_TEMPR41[34] , \R_DATA_TEMPR42[34] , 
        \R_DATA_TEMPR43[34] , \R_DATA_TEMPR44[34] , 
        \R_DATA_TEMPR45[34] , \R_DATA_TEMPR46[34] , 
        \R_DATA_TEMPR47[34] , \R_DATA_TEMPR48[34] , 
        \R_DATA_TEMPR49[34] , \R_DATA_TEMPR50[34] , 
        \R_DATA_TEMPR51[34] , \R_DATA_TEMPR52[34] , 
        \R_DATA_TEMPR53[34] , \R_DATA_TEMPR54[34] , 
        \R_DATA_TEMPR55[34] , \R_DATA_TEMPR56[34] , 
        \R_DATA_TEMPR57[34] , \R_DATA_TEMPR58[34] , 
        \R_DATA_TEMPR59[34] , \R_DATA_TEMPR60[34] , 
        \R_DATA_TEMPR61[34] , \R_DATA_TEMPR62[34] , 
        \R_DATA_TEMPR63[34] , \R_DATA_TEMPR0[35] , \R_DATA_TEMPR1[35] , 
        \R_DATA_TEMPR2[35] , \R_DATA_TEMPR3[35] , \R_DATA_TEMPR4[35] , 
        \R_DATA_TEMPR5[35] , \R_DATA_TEMPR6[35] , \R_DATA_TEMPR7[35] , 
        \R_DATA_TEMPR8[35] , \R_DATA_TEMPR9[35] , \R_DATA_TEMPR10[35] , 
        \R_DATA_TEMPR11[35] , \R_DATA_TEMPR12[35] , 
        \R_DATA_TEMPR13[35] , \R_DATA_TEMPR14[35] , 
        \R_DATA_TEMPR15[35] , \R_DATA_TEMPR16[35] , 
        \R_DATA_TEMPR17[35] , \R_DATA_TEMPR18[35] , 
        \R_DATA_TEMPR19[35] , \R_DATA_TEMPR20[35] , 
        \R_DATA_TEMPR21[35] , \R_DATA_TEMPR22[35] , 
        \R_DATA_TEMPR23[35] , \R_DATA_TEMPR24[35] , 
        \R_DATA_TEMPR25[35] , \R_DATA_TEMPR26[35] , 
        \R_DATA_TEMPR27[35] , \R_DATA_TEMPR28[35] , 
        \R_DATA_TEMPR29[35] , \R_DATA_TEMPR30[35] , 
        \R_DATA_TEMPR31[35] , \R_DATA_TEMPR32[35] , 
        \R_DATA_TEMPR33[35] , \R_DATA_TEMPR34[35] , 
        \R_DATA_TEMPR35[35] , \R_DATA_TEMPR36[35] , 
        \R_DATA_TEMPR37[35] , \R_DATA_TEMPR38[35] , 
        \R_DATA_TEMPR39[35] , \R_DATA_TEMPR40[35] , 
        \R_DATA_TEMPR41[35] , \R_DATA_TEMPR42[35] , 
        \R_DATA_TEMPR43[35] , \R_DATA_TEMPR44[35] , 
        \R_DATA_TEMPR45[35] , \R_DATA_TEMPR46[35] , 
        \R_DATA_TEMPR47[35] , \R_DATA_TEMPR48[35] , 
        \R_DATA_TEMPR49[35] , \R_DATA_TEMPR50[35] , 
        \R_DATA_TEMPR51[35] , \R_DATA_TEMPR52[35] , 
        \R_DATA_TEMPR53[35] , \R_DATA_TEMPR54[35] , 
        \R_DATA_TEMPR55[35] , \R_DATA_TEMPR56[35] , 
        \R_DATA_TEMPR57[35] , \R_DATA_TEMPR58[35] , 
        \R_DATA_TEMPR59[35] , \R_DATA_TEMPR60[35] , 
        \R_DATA_TEMPR61[35] , \R_DATA_TEMPR62[35] , 
        \R_DATA_TEMPR63[35] , \R_DATA_TEMPR0[36] , \R_DATA_TEMPR1[36] , 
        \R_DATA_TEMPR2[36] , \R_DATA_TEMPR3[36] , \R_DATA_TEMPR4[36] , 
        \R_DATA_TEMPR5[36] , \R_DATA_TEMPR6[36] , \R_DATA_TEMPR7[36] , 
        \R_DATA_TEMPR8[36] , \R_DATA_TEMPR9[36] , \R_DATA_TEMPR10[36] , 
        \R_DATA_TEMPR11[36] , \R_DATA_TEMPR12[36] , 
        \R_DATA_TEMPR13[36] , \R_DATA_TEMPR14[36] , 
        \R_DATA_TEMPR15[36] , \R_DATA_TEMPR16[36] , 
        \R_DATA_TEMPR17[36] , \R_DATA_TEMPR18[36] , 
        \R_DATA_TEMPR19[36] , \R_DATA_TEMPR20[36] , 
        \R_DATA_TEMPR21[36] , \R_DATA_TEMPR22[36] , 
        \R_DATA_TEMPR23[36] , \R_DATA_TEMPR24[36] , 
        \R_DATA_TEMPR25[36] , \R_DATA_TEMPR26[36] , 
        \R_DATA_TEMPR27[36] , \R_DATA_TEMPR28[36] , 
        \R_DATA_TEMPR29[36] , \R_DATA_TEMPR30[36] , 
        \R_DATA_TEMPR31[36] , \R_DATA_TEMPR32[36] , 
        \R_DATA_TEMPR33[36] , \R_DATA_TEMPR34[36] , 
        \R_DATA_TEMPR35[36] , \R_DATA_TEMPR36[36] , 
        \R_DATA_TEMPR37[36] , \R_DATA_TEMPR38[36] , 
        \R_DATA_TEMPR39[36] , \R_DATA_TEMPR40[36] , 
        \R_DATA_TEMPR41[36] , \R_DATA_TEMPR42[36] , 
        \R_DATA_TEMPR43[36] , \R_DATA_TEMPR44[36] , 
        \R_DATA_TEMPR45[36] , \R_DATA_TEMPR46[36] , 
        \R_DATA_TEMPR47[36] , \R_DATA_TEMPR48[36] , 
        \R_DATA_TEMPR49[36] , \R_DATA_TEMPR50[36] , 
        \R_DATA_TEMPR51[36] , \R_DATA_TEMPR52[36] , 
        \R_DATA_TEMPR53[36] , \R_DATA_TEMPR54[36] , 
        \R_DATA_TEMPR55[36] , \R_DATA_TEMPR56[36] , 
        \R_DATA_TEMPR57[36] , \R_DATA_TEMPR58[36] , 
        \R_DATA_TEMPR59[36] , \R_DATA_TEMPR60[36] , 
        \R_DATA_TEMPR61[36] , \R_DATA_TEMPR62[36] , 
        \R_DATA_TEMPR63[36] , \R_DATA_TEMPR0[37] , \R_DATA_TEMPR1[37] , 
        \R_DATA_TEMPR2[37] , \R_DATA_TEMPR3[37] , \R_DATA_TEMPR4[37] , 
        \R_DATA_TEMPR5[37] , \R_DATA_TEMPR6[37] , \R_DATA_TEMPR7[37] , 
        \R_DATA_TEMPR8[37] , \R_DATA_TEMPR9[37] , \R_DATA_TEMPR10[37] , 
        \R_DATA_TEMPR11[37] , \R_DATA_TEMPR12[37] , 
        \R_DATA_TEMPR13[37] , \R_DATA_TEMPR14[37] , 
        \R_DATA_TEMPR15[37] , \R_DATA_TEMPR16[37] , 
        \R_DATA_TEMPR17[37] , \R_DATA_TEMPR18[37] , 
        \R_DATA_TEMPR19[37] , \R_DATA_TEMPR20[37] , 
        \R_DATA_TEMPR21[37] , \R_DATA_TEMPR22[37] , 
        \R_DATA_TEMPR23[37] , \R_DATA_TEMPR24[37] , 
        \R_DATA_TEMPR25[37] , \R_DATA_TEMPR26[37] , 
        \R_DATA_TEMPR27[37] , \R_DATA_TEMPR28[37] , 
        \R_DATA_TEMPR29[37] , \R_DATA_TEMPR30[37] , 
        \R_DATA_TEMPR31[37] , \R_DATA_TEMPR32[37] , 
        \R_DATA_TEMPR33[37] , \R_DATA_TEMPR34[37] , 
        \R_DATA_TEMPR35[37] , \R_DATA_TEMPR36[37] , 
        \R_DATA_TEMPR37[37] , \R_DATA_TEMPR38[37] , 
        \R_DATA_TEMPR39[37] , \R_DATA_TEMPR40[37] , 
        \R_DATA_TEMPR41[37] , \R_DATA_TEMPR42[37] , 
        \R_DATA_TEMPR43[37] , \R_DATA_TEMPR44[37] , 
        \R_DATA_TEMPR45[37] , \R_DATA_TEMPR46[37] , 
        \R_DATA_TEMPR47[37] , \R_DATA_TEMPR48[37] , 
        \R_DATA_TEMPR49[37] , \R_DATA_TEMPR50[37] , 
        \R_DATA_TEMPR51[37] , \R_DATA_TEMPR52[37] , 
        \R_DATA_TEMPR53[37] , \R_DATA_TEMPR54[37] , 
        \R_DATA_TEMPR55[37] , \R_DATA_TEMPR56[37] , 
        \R_DATA_TEMPR57[37] , \R_DATA_TEMPR58[37] , 
        \R_DATA_TEMPR59[37] , \R_DATA_TEMPR60[37] , 
        \R_DATA_TEMPR61[37] , \R_DATA_TEMPR62[37] , 
        \R_DATA_TEMPR63[37] , \R_DATA_TEMPR0[38] , \R_DATA_TEMPR1[38] , 
        \R_DATA_TEMPR2[38] , \R_DATA_TEMPR3[38] , \R_DATA_TEMPR4[38] , 
        \R_DATA_TEMPR5[38] , \R_DATA_TEMPR6[38] , \R_DATA_TEMPR7[38] , 
        \R_DATA_TEMPR8[38] , \R_DATA_TEMPR9[38] , \R_DATA_TEMPR10[38] , 
        \R_DATA_TEMPR11[38] , \R_DATA_TEMPR12[38] , 
        \R_DATA_TEMPR13[38] , \R_DATA_TEMPR14[38] , 
        \R_DATA_TEMPR15[38] , \R_DATA_TEMPR16[38] , 
        \R_DATA_TEMPR17[38] , \R_DATA_TEMPR18[38] , 
        \R_DATA_TEMPR19[38] , \R_DATA_TEMPR20[38] , 
        \R_DATA_TEMPR21[38] , \R_DATA_TEMPR22[38] , 
        \R_DATA_TEMPR23[38] , \R_DATA_TEMPR24[38] , 
        \R_DATA_TEMPR25[38] , \R_DATA_TEMPR26[38] , 
        \R_DATA_TEMPR27[38] , \R_DATA_TEMPR28[38] , 
        \R_DATA_TEMPR29[38] , \R_DATA_TEMPR30[38] , 
        \R_DATA_TEMPR31[38] , \R_DATA_TEMPR32[38] , 
        \R_DATA_TEMPR33[38] , \R_DATA_TEMPR34[38] , 
        \R_DATA_TEMPR35[38] , \R_DATA_TEMPR36[38] , 
        \R_DATA_TEMPR37[38] , \R_DATA_TEMPR38[38] , 
        \R_DATA_TEMPR39[38] , \R_DATA_TEMPR40[38] , 
        \R_DATA_TEMPR41[38] , \R_DATA_TEMPR42[38] , 
        \R_DATA_TEMPR43[38] , \R_DATA_TEMPR44[38] , 
        \R_DATA_TEMPR45[38] , \R_DATA_TEMPR46[38] , 
        \R_DATA_TEMPR47[38] , \R_DATA_TEMPR48[38] , 
        \R_DATA_TEMPR49[38] , \R_DATA_TEMPR50[38] , 
        \R_DATA_TEMPR51[38] , \R_DATA_TEMPR52[38] , 
        \R_DATA_TEMPR53[38] , \R_DATA_TEMPR54[38] , 
        \R_DATA_TEMPR55[38] , \R_DATA_TEMPR56[38] , 
        \R_DATA_TEMPR57[38] , \R_DATA_TEMPR58[38] , 
        \R_DATA_TEMPR59[38] , \R_DATA_TEMPR60[38] , 
        \R_DATA_TEMPR61[38] , \R_DATA_TEMPR62[38] , 
        \R_DATA_TEMPR63[38] , \R_DATA_TEMPR0[39] , \R_DATA_TEMPR1[39] , 
        \R_DATA_TEMPR2[39] , \R_DATA_TEMPR3[39] , \R_DATA_TEMPR4[39] , 
        \R_DATA_TEMPR5[39] , \R_DATA_TEMPR6[39] , \R_DATA_TEMPR7[39] , 
        \R_DATA_TEMPR8[39] , \R_DATA_TEMPR9[39] , \R_DATA_TEMPR10[39] , 
        \R_DATA_TEMPR11[39] , \R_DATA_TEMPR12[39] , 
        \R_DATA_TEMPR13[39] , \R_DATA_TEMPR14[39] , 
        \R_DATA_TEMPR15[39] , \R_DATA_TEMPR16[39] , 
        \R_DATA_TEMPR17[39] , \R_DATA_TEMPR18[39] , 
        \R_DATA_TEMPR19[39] , \R_DATA_TEMPR20[39] , 
        \R_DATA_TEMPR21[39] , \R_DATA_TEMPR22[39] , 
        \R_DATA_TEMPR23[39] , \R_DATA_TEMPR24[39] , 
        \R_DATA_TEMPR25[39] , \R_DATA_TEMPR26[39] , 
        \R_DATA_TEMPR27[39] , \R_DATA_TEMPR28[39] , 
        \R_DATA_TEMPR29[39] , \R_DATA_TEMPR30[39] , 
        \R_DATA_TEMPR31[39] , \R_DATA_TEMPR32[39] , 
        \R_DATA_TEMPR33[39] , \R_DATA_TEMPR34[39] , 
        \R_DATA_TEMPR35[39] , \R_DATA_TEMPR36[39] , 
        \R_DATA_TEMPR37[39] , \R_DATA_TEMPR38[39] , 
        \R_DATA_TEMPR39[39] , \R_DATA_TEMPR40[39] , 
        \R_DATA_TEMPR41[39] , \R_DATA_TEMPR42[39] , 
        \R_DATA_TEMPR43[39] , \R_DATA_TEMPR44[39] , 
        \R_DATA_TEMPR45[39] , \R_DATA_TEMPR46[39] , 
        \R_DATA_TEMPR47[39] , \R_DATA_TEMPR48[39] , 
        \R_DATA_TEMPR49[39] , \R_DATA_TEMPR50[39] , 
        \R_DATA_TEMPR51[39] , \R_DATA_TEMPR52[39] , 
        \R_DATA_TEMPR53[39] , \R_DATA_TEMPR54[39] , 
        \R_DATA_TEMPR55[39] , \R_DATA_TEMPR56[39] , 
        \R_DATA_TEMPR57[39] , \R_DATA_TEMPR58[39] , 
        \R_DATA_TEMPR59[39] , \R_DATA_TEMPR60[39] , 
        \R_DATA_TEMPR61[39] , \R_DATA_TEMPR62[39] , 
        \R_DATA_TEMPR63[39] , \BLKX0[0] , \BLKY0[0] , \BLKX1[0] , 
        \BLKY1[0] , \BLKX2[0] , \BLKX2[1] , \BLKX2[2] , \BLKX2[3] , 
        \BLKX2[4] , \BLKX2[5] , \BLKX2[6] , \BLKX2[7] , \BLKX2[8] , 
        \BLKX2[9] , \BLKX2[10] , \BLKX2[11] , \BLKX2[12] , \BLKX2[13] , 
        \BLKX2[14] , \BLKX2[15] , \BLKY2[0] , \BLKY2[1] , \BLKY2[2] , 
        \BLKY2[3] , \BLKY2[4] , \BLKY2[5] , \BLKY2[6] , \BLKY2[7] , 
        \BLKY2[8] , \BLKY2[9] , \BLKY2[10] , \BLKY2[11] , \BLKY2[12] , 
        \BLKY2[13] , \BLKY2[14] , \BLKY2[15] , \ACCESS_BUSY[0][0] , 
        \ACCESS_BUSY[1][0] , \ACCESS_BUSY[2][0] , \ACCESS_BUSY[3][0] , 
        \ACCESS_BUSY[4][0] , \ACCESS_BUSY[5][0] , \ACCESS_BUSY[6][0] , 
        \ACCESS_BUSY[7][0] , \ACCESS_BUSY[8][0] , \ACCESS_BUSY[9][0] , 
        \ACCESS_BUSY[10][0] , \ACCESS_BUSY[11][0] , 
        \ACCESS_BUSY[12][0] , \ACCESS_BUSY[13][0] , 
        \ACCESS_BUSY[14][0] , \ACCESS_BUSY[15][0] , 
        \ACCESS_BUSY[16][0] , \ACCESS_BUSY[17][0] , 
        \ACCESS_BUSY[18][0] , \ACCESS_BUSY[19][0] , 
        \ACCESS_BUSY[20][0] , \ACCESS_BUSY[21][0] , 
        \ACCESS_BUSY[22][0] , \ACCESS_BUSY[23][0] , 
        \ACCESS_BUSY[24][0] , \ACCESS_BUSY[25][0] , 
        \ACCESS_BUSY[26][0] , \ACCESS_BUSY[27][0] , 
        \ACCESS_BUSY[28][0] , \ACCESS_BUSY[29][0] , 
        \ACCESS_BUSY[30][0] , \ACCESS_BUSY[31][0] , 
        \ACCESS_BUSY[32][0] , \ACCESS_BUSY[33][0] , 
        \ACCESS_BUSY[34][0] , \ACCESS_BUSY[35][0] , 
        \ACCESS_BUSY[36][0] , \ACCESS_BUSY[37][0] , 
        \ACCESS_BUSY[38][0] , \ACCESS_BUSY[39][0] , 
        \ACCESS_BUSY[40][0] , \ACCESS_BUSY[41][0] , 
        \ACCESS_BUSY[42][0] , \ACCESS_BUSY[43][0] , 
        \ACCESS_BUSY[44][0] , \ACCESS_BUSY[45][0] , 
        \ACCESS_BUSY[46][0] , \ACCESS_BUSY[47][0] , 
        \ACCESS_BUSY[48][0] , \ACCESS_BUSY[49][0] , 
        \ACCESS_BUSY[50][0] , \ACCESS_BUSY[51][0] , 
        \ACCESS_BUSY[52][0] , \ACCESS_BUSY[53][0] , 
        \ACCESS_BUSY[54][0] , \ACCESS_BUSY[55][0] , 
        \ACCESS_BUSY[56][0] , \ACCESS_BUSY[57][0] , 
        \ACCESS_BUSY[58][0] , \ACCESS_BUSY[59][0] , 
        \ACCESS_BUSY[60][0] , \ACCESS_BUSY[61][0] , 
        \ACCESS_BUSY[62][0] , \ACCESS_BUSY[63][0] , OR4_141_Y, 
        OR4_667_Y, OR4_268_Y, OR4_603_Y, OR4_14_Y, OR4_181_Y, 
        OR4_280_Y, OR4_51_Y, OR4_68_Y, OR4_351_Y, OR4_339_Y, OR4_180_Y, 
        OR4_389_Y, OR4_309_Y, OR4_7_Y, OR4_276_Y, OR4_21_Y, OR4_574_Y, 
        OR4_605_Y, OR4_61_Y, OR4_731_Y, OR4_696_Y, OR4_710_Y, 
        OR4_459_Y, OR4_209_Y, OR4_342_Y, OR4_340_Y, OR4_471_Y, 
        OR4_126_Y, OR4_547_Y, OR4_13_Y, OR4_521_Y, OR4_642_Y, 
        OR4_115_Y, OR4_503_Y, OR4_637_Y, OR4_387_Y, OR4_272_Y, 
        OR4_116_Y, OR4_506_Y, OR4_618_Y, OR4_152_Y, OR4_270_Y, 
        OR4_346_Y, OR4_92_Y, OR4_245_Y, OR4_97_Y, OR4_513_Y, OR4_54_Y, 
        OR4_632_Y, OR4_89_Y, OR4_314_Y, OR4_792_Y, OR4_130_Y, 
        OR4_671_Y, OR4_296_Y, OR4_679_Y, OR4_1_Y, OR4_95_Y, OR4_176_Y, 
        OR4_512_Y, OR4_485_Y, OR4_377_Y, OR4_18_Y, OR4_658_Y, 
        OR4_330_Y, OR4_494_Y, OR4_93_Y, OR4_148_Y, OR4_326_Y, 
        OR4_588_Y, OR4_300_Y, OR4_416_Y, OR4_695_Y, OR4_289_Y, 
        OR4_409_Y, OR4_166_Y, OR4_35_Y, OR4_699_Y, OR4_306_Y, 
        OR4_373_Y, OR4_6_Y, OR4_149_Y, OR4_191_Y, OR4_755_Y, OR4_523_Y, 
        OR4_560_Y, OR4_706_Y, OR4_198_Y, OR4_665_Y, OR4_653_Y, 
        OR4_235_Y, OR4_457_Y, OR4_616_Y, OR4_727_Y, OR4_641_Y, 
        OR4_454_Y, OR4_376_Y, OR4_439_Y, OR4_302_Y, OR4_556_Y, 
        OR4_193_Y, OR4_332_Y, OR4_375_Y, OR4_138_Y, OR4_705_Y, 
        OR4_738_Y, OR4_86_Y, OR4_378_Y, OR4_766_Y, OR4_747_Y, 
        OR4_597_Y, OR4_4_Y, OR4_720_Y, OR4_428_Y, OR4_681_Y, OR4_438_Y, 
        OR4_197_Y, OR4_221_Y, OR4_395_Y, OR4_660_Y, OR4_749_Y, 
        OR4_501_Y, OR4_654_Y, OR4_636_Y, OR4_628_Y, OR4_572_Y, 
        OR4_781_Y, OR4_113_Y, OR4_680_Y, OR4_133_Y, OR4_364_Y, 
        OR4_34_Y, OR4_186_Y, OR4_716_Y, OR4_335_Y, OR4_726_Y, OR4_48_Y, 
        OR4_140_Y, OR4_777_Y, OR4_425_Y, OR4_217_Y, OR4_179_Y, 
        OR4_155_Y, OR4_687_Y, OR4_530_Y, OR4_517_Y, OR4_208_Y, 
        OR4_59_Y, OR4_241_Y, OR4_497_Y, OR4_206_Y, OR4_325_Y, 
        OR4_609_Y, OR4_196_Y, OR4_320_Y, OR4_66_Y, OR4_742_Y, 
        OR4_612_Y, OR4_26_Y, OR4_264_Y, OR4_73_Y, OR4_22_Y, OR4_686_Y, 
        OR4_571_Y, OR4_40_Y, OR4_384_Y, OR4_713_Y, OR4_430_Y, 
        OR4_544_Y, OR4_535_Y, OR4_104_Y, OR4_337_Y, OR4_489_Y, 
        OR4_614_Y, OR4_518_Y, OR4_336_Y, OR4_267_Y, OR4_318_Y, 
        OR4_367_Y, OR4_760_Y, OR4_656_Y, OR4_298_Y, OR4_401_Y, 
        OR4_522_Y, OR4_352_Y, OR4_222_Y, OR4_269_Y, OR4_237_Y, 
        OR4_258_Y, OR4_243_Y, OR4_622_Y, OR4_47_Y, OR4_202_Y, 
        OR4_319_Y, OR4_230_Y, OR4_43_Y, OR4_764_Y, OR4_27_Y, OR4_143_Y, 
        OR4_633_Y, OR4_216_Y, OR4_524_Y, OR4_301_Y, OR4_142_Y, 
        OR4_611_Y, OR4_646_Y, OR4_256_Y, OR4_700_Y, OR4_445_Y, 
        OR4_708_Y, OR4_412_Y, OR4_536_Y, OR4_12_Y, OR4_400_Y, 
        OR4_529_Y, OR4_291_Y, OR4_154_Y, OR4_15_Y, OR4_25_Y, OR4_692_Y, 
        OR4_417_Y, OR4_5_Y, OR4_356_Y, OR4_561_Y, OR4_730_Y, OR4_19_Y, 
        OR4_607_Y, OR4_629_Y, OR4_504_Y, OR4_776_Y, OR4_476_Y, 
        OR4_596_Y, OR4_71_Y, OR4_463_Y, OR4_589_Y, OR4_347_Y, 
        OR4_226_Y, OR4_75_Y, OR4_234_Y, OR4_101_Y, OR4_266_Y, 
        OR4_460_Y, OR4_620_Y, OR4_259_Y, OR4_702_Y, OR4_447_Y, 
        OR4_174_Y, OR4_418_Y, OR4_119_Y, OR4_385_Y, OR4_613_Y, 
        OR4_290_Y, OR4_435_Y, OR4_164_Y, OR4_579_Y, OR4_175_Y, 
        OR4_304_Y, OR4_386_Y, OR4_282_Y, OR4_655_Y, OR4_33_Y, 
        OR4_398_Y, OR4_88_Y, OR4_592_Y, OR4_424_Y, OR4_600_Y, 
        OR4_163_Y, OR4_153_Y, OR4_139_Y, OR4_124_Y, OR4_514_Y, 
        OR4_734_Y, OR4_91_Y, OR4_214_Y, OR4_107_Y, OR4_732_Y, 
        OR4_657_Y, OR4_719_Y, OR4_327_Y, OR4_194_Y, OR4_415_Y, 
        OR4_354_Y, OR4_413_Y, OR4_244_Y, OR4_502_Y, OR4_703_Y, 
        OR4_277_Y, OR4_328_Y, OR4_212_Y, OR4_470_Y, OR4_690_Y, 
        OR4_366_Y, OR4_520_Y, OR4_254_Y, OR4_670_Y, OR4_271_Y, 
        OR4_382_Y, OR4_474_Y, OR4_434_Y, OR4_442_Y, OR4_273_Y, 
        OR4_210_Y, OR4_60_Y, OR4_756_Y, OR4_232_Y, OR4_567_Y, OR4_96_Y, 
        OR4_617_Y, OR4_649_Y, OR4_638_Y, OR4_479_Y, OR4_685_Y, 
        OR4_601_Y, OR4_307_Y, OR4_558_Y, OR4_315_Y, OR4_63_Y, OR4_98_Y, 
        OR4_468_Y, OR4_144_Y, OR4_37_Y, OR4_472_Y, OR4_582_Y, 
        OR4_701_Y, OR4_539_Y, OR4_404_Y, OR4_443_Y, OR4_420_Y, 
        OR4_353_Y, OR4_341_Y, OR4_182_Y, OR4_391_Y, OR4_311_Y, OR4_8_Y, 
        OR4_278_Y, OR4_24_Y, OR4_577_Y, OR4_608_Y, OR4_253_Y, OR4_36_Y, 
        OR4_224_Y, OR4_581_Y, OR4_285_Y, OR4_783_Y, OR4_606_Y, 
        OR4_791_Y, OR4_344_Y, OR4_338_Y, OR4_252_Y, OR4_239_Y, 
        OR4_70_Y, OR4_294_Y, OR4_203_Y, OR4_707_Y, OR4_161_Y, 
        OR4_718_Y, OR4_473_Y, OR4_496_Y, OR4_429_Y, OR4_310_Y, 
        OR4_736_Y, OR4_77_Y, OR4_117_Y, OR4_691_Y, OR4_451_Y, 
        OR4_495_Y, OR4_643_Y, OR4_120_Y, OR4_111_Y, OR4_383_Y, 
        OR4_83_Y, OR4_211_Y, OR4_488_Y, OR4_67_Y, OR4_205_Y, OR4_758_Y, 
        OR4_639_Y, OR4_491_Y, OR4_551_Y, OR4_187_Y, OR4_565_Y, 
        OR4_30_Y, OR4_134_Y, OR4_103_Y, OR4_369_Y, OR4_195_Y, 
        OR4_192_Y, OR4_157_Y, OR4_207_Y, OR4_466_Y, OR4_688_Y, 
        OR4_362_Y, OR4_511_Y, OR4_249_Y, OR4_663_Y, OR4_261_Y, 
        OR4_379_Y, OR4_469_Y, OR4_584_Y, OR4_441_Y, OR4_397_Y, 
        OR4_549_Y, OR4_610_Y, OR4_526_Y, OR4_251_Y, OR4_531_Y, 
        OR4_225_Y, OR4_540_Y, OR4_450_Y, OR4_717_Y, OR4_132_Y, 
        OR4_619_Y, OR4_763_Y, OR4_490_Y, OR4_105_Y, OR4_500_Y, 
        OR4_630_Y, OR4_721_Y, OR4_419_Y, OR4_402_Y, OR4_492_Y, 
        OR4_303_Y, OR4_599_Y, OR4_114_Y, OR4_167_Y, OR4_431_Y, 
        OR4_160_Y, OR4_532_Y, OR4_421_Y, OR4_682_Y, OR4_99_Y, 
        OR4_570_Y, OR4_724_Y, OR4_455_Y, OR4_64_Y, OR4_465_Y, 
        OR4_593_Y, OR4_684_Y, OR4_510_Y, OR4_170_Y, OR4_552_Y, 
        OR4_752_Y, OR4_31_Y, OR4_240_Y, OR4_678_Y, OR4_185_Y, 
        OR4_562_Y, OR4_444_Y, OR4_458_Y, OR4_448_Y, OR4_29_Y, 
        OR4_265_Y, OR4_406_Y, OR4_528_Y, OR4_433_Y, OR4_260_Y, 
        OR4_172_Y, OR4_238_Y, OR4_42_Y, OR4_189_Y, OR4_9_Y, OR4_751_Y, 
        OR4_623_Y, OR4_508_Y, OR4_784_Y, OR4_322_Y, OR4_650_Y, 
        OR4_361_Y, OR4_797_Y, OR4_274_Y, OR4_773_Y, OR4_85_Y, 
        OR4_371_Y, OR4_750_Y, OR4_78_Y, OR4_645_Y, OR4_515_Y, 
        OR4_372_Y, OR4_626_Y, OR4_694_Y, OR4_587_Y, OR4_229_Y, 
        OR4_334_Y, OR4_449_Y, OR4_292_Y, OR4_151_Y, OR4_190_Y, 
        OR4_165_Y, OR4_505_Y, OR4_779_Y, OR4_477_Y, OR4_598_Y, 
        OR4_72_Y, OR4_464_Y, OR4_591_Y, OR4_350_Y, OR4_227_Y, OR4_76_Y, 
        OR4_405_Y, OR4_585_Y, OR4_774_Y, OR4_331_Y, OR4_28_Y, 
        OR4_527_Y, OR4_358_Y, OR4_537_Y, OR4_94_Y, OR4_87_Y, OR4_403_Y, 
        OR4_669_Y, OR4_368_Y, OR4_487_Y, OR4_780_Y, OR4_359_Y, 
        OR4_481_Y, OR4_250_Y, OR4_106_Y, OR4_782_Y, OR4_580_Y, OR4_0_Y, 
        OR4_765_Y, OR4_785_Y, OR4_534_Y, OR4_283_Y, OR4_410_Y, 
        OR4_408_Y, OR4_541_Y, OR4_201_Y, OR4_299_Y, OR4_286_Y, 
        OR4_662_Y, OR4_84_Y, OR4_246_Y, OR4_360_Y, OR4_275_Y, OR4_81_Y, 
        OR4_3_Y, OR4_56_Y, OR4_263_Y, OR4_123_Y, OR4_759_Y, OR4_507_Y, 
        OR4_664_Y, OR4_365_Y, OR4_640_Y, OR4_566_Y, OR4_247_Y, 
        OR4_121_Y, OR4_147_Y, OR4_411_Y, OR4_634_Y, OR4_308_Y, 
        OR4_452_Y, OR4_183_Y, OR4_604_Y, OR4_199_Y, OR4_323_Y, 
        OR4_414_Y, OR4_789_Y, OR4_357_Y, OR4_733_Y, OR4_135_Y, 
        OR4_218_Y, OR4_422_Y, OR4_53_Y, OR4_370_Y, OR4_745_Y, 
        OR4_625_Y, OR4_557_Y, OR4_546_Y, OR4_388_Y, OR4_602_Y, 
        OR4_516_Y, OR4_223_Y, OR4_475_Y, OR4_236_Y, OR4_793_Y, 
        OR4_10_Y, OR4_137_Y, OR4_573_Y, OR4_554_Y, OR4_446_Y, OR4_80_Y, 
        OR4_723_Y, OR4_394_Y, OR4_559_Y, OR4_162_Y, OR4_219_Y, 
        OR4_58_Y, OR4_49_Y, OR4_440_Y, OR4_666_Y, OR4_16_Y, OR4_128_Y, 
        OR4_39_Y, OR4_661_Y, OR4_575_Y, OR4_647_Y, OR4_46_Y, OR4_188_Y, 
        OR4_146_Y, OR4_159_Y, OR4_712_Y, OR4_456_Y, OR4_594_Y, 
        OR4_590_Y, OR4_722_Y, OR4_380_Y, OR4_390_Y, OR4_381_Y, 
        OR4_233_Y, OR4_437_Y, OR4_348_Y, OR4_50_Y, OR4_313_Y, OR4_55_Y, 
        OR4_624_Y, OR4_651_Y, OR4_355_Y, CFG3_10_Y, CFG3_9_Y, CFG3_0_Y, 
        CFG3_12_Y, CFG3_11_Y, CFG3_6_Y, CFG3_1_Y, CFG3_13_Y, CFG2_0_Y, 
        CFG2_1_Y, OR4_762_Y, OR4_735_Y, OR4_627_Y, OR4_279_Y, 
        OR4_102_Y, OR4_576_Y, OR4_737_Y, OR4_343_Y, OR4_399_Y, 
        OR4_169_Y, OR4_158_Y, OR4_799_Y, OR4_213_Y, OR4_118_Y, 
        OR4_631_Y, OR4_79_Y, OR4_644_Y, OR4_396_Y, OR4_427_Y, 
        OR4_145_Y, OR4_484_Y, OR4_288_Y, OR4_255_Y, OR4_231_Y, 
        OR4_748_Y, OR4_595_Y, OR4_578_Y, OR4_281_Y, OR4_129_Y, 
        OR4_787_Y, OR4_767_Y, OR4_345_Y, OR4_569_Y, OR4_725_Y, 
        OR4_44_Y, OR4_744_Y, OR4_568_Y, OR4_486_Y, OR4_550_Y, 
        OR4_564_Y, OR4_467_Y, OR4_728_Y, OR4_509_Y, OR4_392_Y, 
        OR4_772_Y, OR4_108_Y, OR4_583_Y, OR4_493_Y, OR4_220_Y, 
        OR4_482_Y, OR4_741_Y, OR4_171_Y, OR4_648_Y, OR4_794_Y, 
        OR4_525_Y, OR4_136_Y, OR4_538_Y, OR4_659_Y, OR4_746_Y, 
        OR4_740_Y, OR4_697_Y, OR4_287_Y, OR4_586_Y, OR4_363_Y, 
        OR4_215_Y, OR4_677_Y, OR4_709_Y, OR4_316_Y, OR4_771_Y, 
        OR4_184_Y, OR4_173_Y, OR4_553_Y, OR4_790_Y, OR4_127_Y, 
        OR4_262_Y, OR4_156_Y, OR4_788_Y, OR4_698_Y, OR4_754_Y, 
        OR4_563_Y, OR4_757_Y, OR4_480_Y, OR4_62_Y, OR4_423_Y, 
        OR4_635_Y, OR4_798_Y, OR4_82_Y, OR4_674_Y, OR4_693_Y, 
        OR4_257_Y, OR4_242_Y, OR4_621_Y, OR4_45_Y, OR4_200_Y, 
        OR4_317_Y, OR4_228_Y, OR4_41_Y, OR4_761_Y, OR4_23_Y, OR4_775_Y, 
        CFG3_7_Y, CFG3_4_Y, CFG3_8_Y, CFG3_2_Y, CFG3_3_Y, CFG3_14_Y, 
        CFG3_5_Y, CFG3_15_Y, CFG2_2_Y, CFG2_3_Y, OR4_100_Y, OR4_483_Y, 
        OR4_689_Y, OR4_768_Y, OR4_168_Y, OR4_615_Y, OR4_110_Y, 
        OR4_499_Y, OR4_374_Y, OR4_715_Y, OR4_178_Y, OR4_683_Y, OR4_2_Y, 
        OR4_295_Y, OR4_676_Y, OR4_796_Y, OR4_555_Y, OR4_432_Y, 
        OR4_297_Y, OR4_305_Y, OR4_652_Y, OR4_743_Y, OR4_533_Y, 
        OR4_426_Y, OR4_729_Y, OR4_11_Y, OR4_65_Y, OR4_17_Y, OR4_478_Y, 
        OR4_668_Y, OR4_122_Y, OR4_349_Y, OR4_20_Y, OR4_177_Y, 
        OR4_704_Y, OR4_324_Y, OR4_714_Y, OR4_38_Y, OR4_125_Y, 
        OR4_770_Y, OR4_675_Y, OR4_462_Y, OR4_436_Y, OR4_407_Y, 
        OR4_131_Y, OR4_786_Y, OR4_769_Y, OR4_453_Y, OR4_321_Y, 
        OR4_69_Y, OR4_57_Y, OR4_711_Y, OR4_112_Y, OR4_32_Y, OR4_542_Y, 
        OR4_795_Y, OR4_548_Y, OR4_312_Y, OR4_333_Y, OR4_673_Y, 
        OR4_74_Y, OR4_461_Y, OR4_778_Y, OR4_545_Y, OR4_393_Y, OR4_52_Y, 
        OR4_90_Y, OR4_498_Y, OR4_150_Y, OR4_293_Y, OR4_284_Y, 
        OR4_109_Y, OR4_329_Y, OR4_248_Y, OR4_739_Y, OR4_204_Y, 
        OR4_753_Y, OR4_519_Y, OR4_543_Y, OR4_672_Y, VCC, GND, 
        ADLIB_VCC;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    assign ADLIB_VCC = VCC_power_net1;
    
    OR4 OR4_700 (.A(\R_DATA_TEMPR16[25] ), .B(\R_DATA_TEMPR17[25] ), 
        .C(\R_DATA_TEMPR18[25] ), .D(\R_DATA_TEMPR19[25] ), .Y(
        OR4_700_Y));
    OR4 OR4_399 (.A(\R_DATA_TEMPR16[32] ), .B(\R_DATA_TEMPR17[32] ), 
        .C(\R_DATA_TEMPR18[32] ), .D(\R_DATA_TEMPR19[32] ), .Y(
        OR4_399_Y));
    OR4 OR4_420 (.A(\R_DATA_TEMPR16[38] ), .B(\R_DATA_TEMPR17[38] ), 
        .C(\R_DATA_TEMPR18[38] ), .D(\R_DATA_TEMPR19[38] ), .Y(
        OR4_420_Y));
    OR4 OR4_738 (.A(\R_DATA_TEMPR8[36] ), .B(\R_DATA_TEMPR9[36] ), .C(
        \R_DATA_TEMPR10[36] ), .D(\R_DATA_TEMPR11[36] ), .Y(OR4_738_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[1]  (.A(CFG3_9_Y), .B(CFG2_0_Y), 
        .Y(\BLKY2[1] ));
    OR4 OR4_402 (.A(OR4_114_Y), .B(OR4_167_Y), .C(OR4_431_Y), .D(
        OR4_160_Y), .Y(OR4_402_Y));
    OR4 OR4_384 (.A(\R_DATA_TEMPR8[19] ), .B(\R_DATA_TEMPR9[19] ), .C(
        \R_DATA_TEMPR10[19] ), .D(\R_DATA_TEMPR11[19] ), .Y(OR4_384_Y));
    OR4 OR4_373 (.A(OR4_755_Y), .B(OR4_523_Y), .C(OR4_560_Y), .D(
        OR4_706_Y), .Y(OR4_373_Y));
    OR4 OR4_770 (.A(\R_DATA_TEMPR60[1] ), .B(\R_DATA_TEMPR61[1] ), .C(
        \R_DATA_TEMPR62[1] ), .D(\R_DATA_TEMPR63[1] ), .Y(OR4_770_Y));
    OR4 OR4_253 (.A(\R_DATA_TEMPR60[38] ), .B(\R_DATA_TEMPR61[38] ), 
        .C(\R_DATA_TEMPR62[38] ), .D(\R_DATA_TEMPR63[38] ), .Y(
        OR4_253_Y));
    OR4 OR4_409 (.A(\R_DATA_TEMPR44[22] ), .B(\R_DATA_TEMPR45[22] ), 
        .C(\R_DATA_TEMPR46[22] ), .D(\R_DATA_TEMPR47[22] ), .Y(
        OR4_409_Y));
    OR4 OR4_472 (.A(OR4_391_Y), .B(OR4_311_Y), .C(OR4_8_Y), .D(
        OR4_278_Y), .Y(OR4_472_Y));
    OR4 OR4_181 (.A(\R_DATA_TEMPR4[34] ), .B(\R_DATA_TEMPR5[34] ), .C(
        \R_DATA_TEMPR6[34] ), .D(\R_DATA_TEMPR7[34] ), .Y(OR4_181_Y));
    OR4 OR4_106 (.A(\R_DATA_TEMPR52[20] ), .B(\R_DATA_TEMPR53[20] ), 
        .C(\R_DATA_TEMPR54[20] ), .D(\R_DATA_TEMPR55[20] ), .Y(
        OR4_106_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%21%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R21C0 (
        .A_DOUT({\R_DATA_TEMPR21[39] , \R_DATA_TEMPR21[38] , 
        \R_DATA_TEMPR21[37] , \R_DATA_TEMPR21[36] , 
        \R_DATA_TEMPR21[35] , \R_DATA_TEMPR21[34] , 
        \R_DATA_TEMPR21[33] , \R_DATA_TEMPR21[32] , 
        \R_DATA_TEMPR21[31] , \R_DATA_TEMPR21[30] , 
        \R_DATA_TEMPR21[29] , \R_DATA_TEMPR21[28] , 
        \R_DATA_TEMPR21[27] , \R_DATA_TEMPR21[26] , 
        \R_DATA_TEMPR21[25] , \R_DATA_TEMPR21[24] , 
        \R_DATA_TEMPR21[23] , \R_DATA_TEMPR21[22] , 
        \R_DATA_TEMPR21[21] , \R_DATA_TEMPR21[20] }), .B_DOUT({
        \R_DATA_TEMPR21[19] , \R_DATA_TEMPR21[18] , 
        \R_DATA_TEMPR21[17] , \R_DATA_TEMPR21[16] , 
        \R_DATA_TEMPR21[15] , \R_DATA_TEMPR21[14] , 
        \R_DATA_TEMPR21[13] , \R_DATA_TEMPR21[12] , 
        \R_DATA_TEMPR21[11] , \R_DATA_TEMPR21[10] , 
        \R_DATA_TEMPR21[9] , \R_DATA_TEMPR21[8] , \R_DATA_TEMPR21[7] , 
        \R_DATA_TEMPR21[6] , \R_DATA_TEMPR21[5] , \R_DATA_TEMPR21[4] , 
        \R_DATA_TEMPR21[3] , \R_DATA_TEMPR21[2] , \R_DATA_TEMPR21[1] , 
        \R_DATA_TEMPR21[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[5] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_83 (.A(\R_DATA_TEMPR28[26] ), .B(\R_DATA_TEMPR29[26] ), .C(
        \R_DATA_TEMPR30[26] ), .D(\R_DATA_TEMPR31[26] ), .Y(OR4_83_Y));
    OR4 OR4_479 (.A(\R_DATA_TEMPR28[39] ), .B(\R_DATA_TEMPR29[39] ), 
        .C(\R_DATA_TEMPR30[39] ), .D(\R_DATA_TEMPR31[39] ), .Y(
        OR4_479_Y));
    OR4 OR4_138 (.A(\R_DATA_TEMPR0[36] ), .B(\R_DATA_TEMPR1[36] ), .C(
        \R_DATA_TEMPR2[36] ), .D(\R_DATA_TEMPR3[36] ), .Y(OR4_138_Y));
    OR4 OR4_176 (.A(\R_DATA_TEMPR60[4] ), .B(\R_DATA_TEMPR61[4] ), .C(
        \R_DATA_TEMPR62[4] ), .D(\R_DATA_TEMPR63[4] ), .Y(OR4_176_Y));
    OR4 OR4_610 (.A(OR4_500_Y), .B(OR4_630_Y), .C(OR4_721_Y), .D(
        OR4_419_Y), .Y(OR4_610_Y));
    OR4 OR4_481 (.A(\R_DATA_TEMPR44[20] ), .B(\R_DATA_TEMPR45[20] ), 
        .C(\R_DATA_TEMPR46[20] ), .D(\R_DATA_TEMPR47[20] ), .Y(
        OR4_481_Y));
    OR4 OR4_488 (.A(\R_DATA_TEMPR36[26] ), .B(\R_DATA_TEMPR37[26] ), 
        .C(\R_DATA_TEMPR38[26] ), .D(\R_DATA_TEMPR39[26] ), .Y(
        OR4_488_Y));
    OR4 OR4_308 (.A(\R_DATA_TEMPR32[5] ), .B(\R_DATA_TEMPR33[5] ), .C(
        \R_DATA_TEMPR34[5] ), .D(\R_DATA_TEMPR35[5] ), .Y(OR4_308_Y));
    OR4 OR4_317 (.A(\R_DATA_TEMPR40[14] ), .B(\R_DATA_TEMPR41[14] ), 
        .C(\R_DATA_TEMPR42[14] ), .D(\R_DATA_TEMPR43[14] ), .Y(
        OR4_317_Y));
    OR4 OR4_110 (.A(\R_DATA_TEMPR8[27] ), .B(\R_DATA_TEMPR9[27] ), .C(
        \R_DATA_TEMPR10[27] ), .D(\R_DATA_TEMPR11[27] ), .Y(OR4_110_Y));
    OR4 OR4_658 (.A(\R_DATA_TEMPR0[22] ), .B(\R_DATA_TEMPR1[22] ), .C(
        \R_DATA_TEMPR2[22] ), .D(\R_DATA_TEMPR3[22] ), .Y(OR4_658_Y));
    OR4 OR4_799 (.A(\R_DATA_TEMPR28[32] ), .B(\R_DATA_TEMPR29[32] ), 
        .C(\R_DATA_TEMPR30[32] ), .D(\R_DATA_TEMPR31[32] ), .Y(
        OR4_799_Y));
    OR4 OR4_378 (.A(\R_DATA_TEMPR16[36] ), .B(\R_DATA_TEMPR17[36] ), 
        .C(\R_DATA_TEMPR18[36] ), .D(\R_DATA_TEMPR19[36] ), .Y(
        OR4_378_Y));
    OR4 OR4_2 (.A(\R_DATA_TEMPR32[27] ), .B(\R_DATA_TEMPR33[27] ), .C(
        \R_DATA_TEMPR34[27] ), .D(\R_DATA_TEMPR35[27] ), .Y(OR4_2_Y));
    OR4 OR4_718 (.A(\R_DATA_TEMPR48[30] ), .B(\R_DATA_TEMPR49[30] ), 
        .C(\R_DATA_TEMPR50[30] ), .D(\R_DATA_TEMPR51[30] ), .Y(
        OR4_718_Y));
    OR4 OR4_329 (.A(\R_DATA_TEMPR32[35] ), .B(\R_DATA_TEMPR33[35] ), 
        .C(\R_DATA_TEMPR34[35] ), .D(\R_DATA_TEMPR35[35] ), .Y(
        OR4_329_Y));
    OR4 \OR4_R_DATA[29]  (.A(OR4_189_Y), .B(OR4_9_Y), .C(OR4_751_Y), 
        .D(OR4_623_Y), .Y(R_DATA[29]));
    OR4 OR4_765 (.A(OR4_201_Y), .B(OR4_299_Y), .C(OR4_286_Y), .D(
        OR4_662_Y), .Y(OR4_765_Y));
    OR4 OR4_667 (.A(OR4_68_Y), .B(OR4_351_Y), .C(OR4_339_Y), .D(
        OR4_180_Y), .Y(OR4_667_Y));
    OR4 OR4_652 (.A(OR4_729_Y), .B(OR4_11_Y), .C(OR4_65_Y), .D(
        OR4_17_Y), .Y(OR4_652_Y));
    OR4 OR4_766 (.A(\R_DATA_TEMPR20[36] ), .B(\R_DATA_TEMPR21[36] ), 
        .C(\R_DATA_TEMPR22[36] ), .D(\R_DATA_TEMPR23[36] ), .Y(
        OR4_766_Y));
    OR4 OR4_593 (.A(\R_DATA_TEMPR52[8] ), .B(\R_DATA_TEMPR53[8] ), .C(
        \R_DATA_TEMPR54[8] ), .D(\R_DATA_TEMPR55[8] ), .Y(OR4_593_Y));
    OR4 OR4_48 (.A(\R_DATA_TEMPR52[0] ), .B(\R_DATA_TEMPR53[0] ), .C(
        \R_DATA_TEMPR54[0] ), .D(\R_DATA_TEMPR55[0] ), .Y(OR4_48_Y));
    OR4 OR4_589 (.A(\R_DATA_TEMPR44[24] ), .B(\R_DATA_TEMPR45[24] ), 
        .C(\R_DATA_TEMPR46[24] ), .D(\R_DATA_TEMPR47[24] ), .Y(
        OR4_589_Y));
    OR4 OR4_109 (.A(\R_DATA_TEMPR28[35] ), .B(\R_DATA_TEMPR29[35] ), 
        .C(\R_DATA_TEMPR30[35] ), .D(\R_DATA_TEMPR31[35] ), .Y(
        OR4_109_Y));
    OR4 OR4_241 (.A(\R_DATA_TEMPR20[23] ), .B(\R_DATA_TEMPR21[23] ), 
        .C(\R_DATA_TEMPR22[23] ), .D(\R_DATA_TEMPR23[23] ), .Y(
        OR4_241_Y));
    OR4 OR4_580 (.A(\R_DATA_TEMPR60[20] ), .B(\R_DATA_TEMPR61[20] ), 
        .C(\R_DATA_TEMPR62[20] ), .D(\R_DATA_TEMPR63[20] ), .Y(
        OR4_580_Y));
    OR4 OR4_81 (.A(\R_DATA_TEMPR48[11] ), .B(\R_DATA_TEMPR49[11] ), .C(
        \R_DATA_TEMPR50[11] ), .D(\R_DATA_TEMPR51[11] ), .Y(OR4_81_Y));
    OR4 OR4_118 (.A(\R_DATA_TEMPR36[32] ), .B(\R_DATA_TEMPR37[32] ), 
        .C(\R_DATA_TEMPR38[32] ), .D(\R_DATA_TEMPR39[32] ), .Y(
        OR4_118_Y));
    OR4 \OR4_R_DATA[7]  (.A(OR4_467_Y), .B(OR4_728_Y), .C(OR4_509_Y), 
        .D(OR4_392_Y), .Y(R_DATA[7]));
    OR4 OR4_179 (.A(OR4_325_Y), .B(OR4_609_Y), .C(OR4_196_Y), .D(
        OR4_320_Y), .Y(OR4_179_Y));
    OR4 OR4_542 (.A(\R_DATA_TEMPR40[33] ), .B(\R_DATA_TEMPR41[33] ), 
        .C(\R_DATA_TEMPR42[33] ), .D(\R_DATA_TEMPR43[33] ), .Y(
        OR4_542_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R54C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%54%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R54C0 (
        .A_DOUT({\R_DATA_TEMPR54[39] , \R_DATA_TEMPR54[38] , 
        \R_DATA_TEMPR54[37] , \R_DATA_TEMPR54[36] , 
        \R_DATA_TEMPR54[35] , \R_DATA_TEMPR54[34] , 
        \R_DATA_TEMPR54[33] , \R_DATA_TEMPR54[32] , 
        \R_DATA_TEMPR54[31] , \R_DATA_TEMPR54[30] , 
        \R_DATA_TEMPR54[29] , \R_DATA_TEMPR54[28] , 
        \R_DATA_TEMPR54[27] , \R_DATA_TEMPR54[26] , 
        \R_DATA_TEMPR54[25] , \R_DATA_TEMPR54[24] , 
        \R_DATA_TEMPR54[23] , \R_DATA_TEMPR54[22] , 
        \R_DATA_TEMPR54[21] , \R_DATA_TEMPR54[20] }), .B_DOUT({
        \R_DATA_TEMPR54[19] , \R_DATA_TEMPR54[18] , 
        \R_DATA_TEMPR54[17] , \R_DATA_TEMPR54[16] , 
        \R_DATA_TEMPR54[15] , \R_DATA_TEMPR54[14] , 
        \R_DATA_TEMPR54[13] , \R_DATA_TEMPR54[12] , 
        \R_DATA_TEMPR54[11] , \R_DATA_TEMPR54[10] , 
        \R_DATA_TEMPR54[9] , \R_DATA_TEMPR54[8] , \R_DATA_TEMPR54[7] , 
        \R_DATA_TEMPR54[6] , \R_DATA_TEMPR54[5] , \R_DATA_TEMPR54[4] , 
        \R_DATA_TEMPR54[3] , \R_DATA_TEMPR54[2] , \R_DATA_TEMPR54[1] , 
        \R_DATA_TEMPR54[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[54][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[13] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[13] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R45C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%45%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R45C0 (
        .A_DOUT({\R_DATA_TEMPR45[39] , \R_DATA_TEMPR45[38] , 
        \R_DATA_TEMPR45[37] , \R_DATA_TEMPR45[36] , 
        \R_DATA_TEMPR45[35] , \R_DATA_TEMPR45[34] , 
        \R_DATA_TEMPR45[33] , \R_DATA_TEMPR45[32] , 
        \R_DATA_TEMPR45[31] , \R_DATA_TEMPR45[30] , 
        \R_DATA_TEMPR45[29] , \R_DATA_TEMPR45[28] , 
        \R_DATA_TEMPR45[27] , \R_DATA_TEMPR45[26] , 
        \R_DATA_TEMPR45[25] , \R_DATA_TEMPR45[24] , 
        \R_DATA_TEMPR45[23] , \R_DATA_TEMPR45[22] , 
        \R_DATA_TEMPR45[21] , \R_DATA_TEMPR45[20] }), .B_DOUT({
        \R_DATA_TEMPR45[19] , \R_DATA_TEMPR45[18] , 
        \R_DATA_TEMPR45[17] , \R_DATA_TEMPR45[16] , 
        \R_DATA_TEMPR45[15] , \R_DATA_TEMPR45[14] , 
        \R_DATA_TEMPR45[13] , \R_DATA_TEMPR45[12] , 
        \R_DATA_TEMPR45[11] , \R_DATA_TEMPR45[10] , 
        \R_DATA_TEMPR45[9] , \R_DATA_TEMPR45[8] , \R_DATA_TEMPR45[7] , 
        \R_DATA_TEMPR45[6] , \R_DATA_TEMPR45[5] , \R_DATA_TEMPR45[4] , 
        \R_DATA_TEMPR45[3] , \R_DATA_TEMPR45[2] , \R_DATA_TEMPR45[1] , 
        \R_DATA_TEMPR45[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[45][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[11] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[11] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_729 (.A(\R_DATA_TEMPR0[1] ), .B(\R_DATA_TEMPR1[1] ), .C(
        \R_DATA_TEMPR2[1] ), .D(\R_DATA_TEMPR3[1] ), .Y(OR4_729_Y));
    OR4 \OR4_R_DATA[4]  (.A(OR4_618_Y), .B(OR4_152_Y), .C(OR4_270_Y), 
        .D(OR4_346_Y), .Y(R_DATA[4]));
    OR4 OR4_135 (.A(OR4_602_Y), .B(OR4_516_Y), .C(OR4_223_Y), .D(
        OR4_475_Y), .Y(OR4_135_Y));
    OR4 OR4_383 (.A(\R_DATA_TEMPR24[26] ), .B(\R_DATA_TEMPR25[26] ), 
        .C(\R_DATA_TEMPR26[26] ), .D(\R_DATA_TEMPR27[26] ), .Y(
        OR4_383_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[9]  (.A(CFG3_9_Y), .B(CFG2_1_Y), 
        .Y(\BLKY2[9] ));
    OR4 OR4_780 (.A(\R_DATA_TEMPR36[20] ), .B(\R_DATA_TEMPR37[20] ), 
        .C(\R_DATA_TEMPR38[20] ), .D(\R_DATA_TEMPR39[20] ), .Y(
        OR4_780_Y));
    OR4 OR4_544 (.A(\R_DATA_TEMPR20[19] ), .B(\R_DATA_TEMPR21[19] ), 
        .C(\R_DATA_TEMPR22[19] ), .D(\R_DATA_TEMPR23[19] ), .Y(
        OR4_544_Y));
    OR4 OR4_267 (.A(\R_DATA_TEMPR52[19] ), .B(\R_DATA_TEMPR53[19] ), 
        .C(\R_DATA_TEMPR54[19] ), .D(\R_DATA_TEMPR55[19] ), .Y(
        OR4_267_Y));
    CFG3 #( .INIT(8'h10) )  CFG3_9 (.A(R_ADDR[13]), .B(R_ADDR[12]), .C(
        R_ADDR[11]), .Y(CFG3_9_Y));
    OR4 OR4_523 (.A(\R_DATA_TEMPR4[16] ), .B(\R_DATA_TEMPR5[16] ), .C(
        \R_DATA_TEMPR6[16] ), .D(\R_DATA_TEMPR7[16] ), .Y(OR4_523_Y));
    OR4 OR4_437 (.A(\R_DATA_TEMPR32[31] ), .B(\R_DATA_TEMPR33[31] ), 
        .C(\R_DATA_TEMPR34[31] ), .D(\R_DATA_TEMPR35[31] ), .Y(
        OR4_437_Y));
    OR4 OR4_482 (.A(\R_DATA_TEMPR20[7] ), .B(\R_DATA_TEMPR21[7] ), .C(
        \R_DATA_TEMPR22[7] ), .D(\R_DATA_TEMPR23[7] ), .Y(OR4_482_Y));
    OR4 OR4_167 (.A(\R_DATA_TEMPR4[8] ), .B(\R_DATA_TEMPR5[8] ), .C(
        \R_DATA_TEMPR6[8] ), .D(\R_DATA_TEMPR7[8] ), .Y(OR4_167_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R51C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%51%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R51C0 (
        .A_DOUT({\R_DATA_TEMPR51[39] , \R_DATA_TEMPR51[38] , 
        \R_DATA_TEMPR51[37] , \R_DATA_TEMPR51[36] , 
        \R_DATA_TEMPR51[35] , \R_DATA_TEMPR51[34] , 
        \R_DATA_TEMPR51[33] , \R_DATA_TEMPR51[32] , 
        \R_DATA_TEMPR51[31] , \R_DATA_TEMPR51[30] , 
        \R_DATA_TEMPR51[29] , \R_DATA_TEMPR51[28] , 
        \R_DATA_TEMPR51[27] , \R_DATA_TEMPR51[26] , 
        \R_DATA_TEMPR51[25] , \R_DATA_TEMPR51[24] , 
        \R_DATA_TEMPR51[23] , \R_DATA_TEMPR51[22] , 
        \R_DATA_TEMPR51[21] , \R_DATA_TEMPR51[20] }), .B_DOUT({
        \R_DATA_TEMPR51[19] , \R_DATA_TEMPR51[18] , 
        \R_DATA_TEMPR51[17] , \R_DATA_TEMPR51[16] , 
        \R_DATA_TEMPR51[15] , \R_DATA_TEMPR51[14] , 
        \R_DATA_TEMPR51[13] , \R_DATA_TEMPR51[12] , 
        \R_DATA_TEMPR51[11] , \R_DATA_TEMPR51[10] , 
        \R_DATA_TEMPR51[9] , \R_DATA_TEMPR51[8] , \R_DATA_TEMPR51[7] , 
        \R_DATA_TEMPR51[6] , \R_DATA_TEMPR51[5] , \R_DATA_TEMPR51[4] , 
        \R_DATA_TEMPR51[3] , \R_DATA_TEMPR51[2] , \R_DATA_TEMPR51[1] , 
        \R_DATA_TEMPR51[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[51][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[12] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[12] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_705 (.A(\R_DATA_TEMPR4[36] ), .B(\R_DATA_TEMPR5[36] ), .C(
        \R_DATA_TEMPR6[36] ), .D(\R_DATA_TEMPR7[36] ), .Y(OR4_705_Y));
    OR4 OR4_607 (.A(\R_DATA_TEMPR12[24] ), .B(\R_DATA_TEMPR13[24] ), 
        .C(\R_DATA_TEMPR14[24] ), .D(\R_DATA_TEMPR15[24] ), .Y(
        OR4_607_Y));
    OR4 OR4_489 (.A(\R_DATA_TEMPR36[19] ), .B(\R_DATA_TEMPR37[19] ), 
        .C(\R_DATA_TEMPR38[19] ), .D(\R_DATA_TEMPR39[19] ), .Y(
        OR4_489_Y));
    OR4 OR4_706 (.A(\R_DATA_TEMPR12[16] ), .B(\R_DATA_TEMPR13[16] ), 
        .C(\R_DATA_TEMPR14[16] ), .D(\R_DATA_TEMPR15[16] ), .Y(
        OR4_706_Y));
    OR4 OR4_186 (.A(\R_DATA_TEMPR36[0] ), .B(\R_DATA_TEMPR37[0] ), .C(
        \R_DATA_TEMPR38[0] ), .D(\R_DATA_TEMPR39[0] ), .Y(OR4_186_Y));
    OR4 OR4_775 (.A(\R_DATA_TEMPR60[14] ), .B(\R_DATA_TEMPR61[14] ), 
        .C(\R_DATA_TEMPR62[14] ), .D(\R_DATA_TEMPR63[14] ), .Y(
        OR4_775_Y));
    OR4 OR4_677 (.A(\R_DATA_TEMPR4[15] ), .B(\R_DATA_TEMPR5[15] ), .C(
        \R_DATA_TEMPR6[15] ), .D(\R_DATA_TEMPR7[15] ), .Y(OR4_677_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%6%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R6C0 (.A_DOUT({
        \R_DATA_TEMPR6[39] , \R_DATA_TEMPR6[38] , \R_DATA_TEMPR6[37] , 
        \R_DATA_TEMPR6[36] , \R_DATA_TEMPR6[35] , \R_DATA_TEMPR6[34] , 
        \R_DATA_TEMPR6[33] , \R_DATA_TEMPR6[32] , \R_DATA_TEMPR6[31] , 
        \R_DATA_TEMPR6[30] , \R_DATA_TEMPR6[29] , \R_DATA_TEMPR6[28] , 
        \R_DATA_TEMPR6[27] , \R_DATA_TEMPR6[26] , \R_DATA_TEMPR6[25] , 
        \R_DATA_TEMPR6[24] , \R_DATA_TEMPR6[23] , \R_DATA_TEMPR6[22] , 
        \R_DATA_TEMPR6[21] , \R_DATA_TEMPR6[20] }), .B_DOUT({
        \R_DATA_TEMPR6[19] , \R_DATA_TEMPR6[18] , \R_DATA_TEMPR6[17] , 
        \R_DATA_TEMPR6[16] , \R_DATA_TEMPR6[15] , \R_DATA_TEMPR6[14] , 
        \R_DATA_TEMPR6[13] , \R_DATA_TEMPR6[12] , \R_DATA_TEMPR6[11] , 
        \R_DATA_TEMPR6[10] , \R_DATA_TEMPR6[9] , \R_DATA_TEMPR6[8] , 
        \R_DATA_TEMPR6[7] , \R_DATA_TEMPR6[6] , \R_DATA_TEMPR6[5] , 
        \R_DATA_TEMPR6[4] , \R_DATA_TEMPR6[3] , \R_DATA_TEMPR6[2] , 
        \R_DATA_TEMPR6[1] , \R_DATA_TEMPR6[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[6][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_235 (.A(\R_DATA_TEMPR28[16] ), .B(\R_DATA_TEMPR29[16] ), 
        .C(\R_DATA_TEMPR30[16] ), .D(\R_DATA_TEMPR31[16] ), .Y(
        OR4_235_Y));
    OR4 OR4_341 (.A(\R_DATA_TEMPR24[38] ), .B(\R_DATA_TEMPR25[38] ), 
        .C(\R_DATA_TEMPR26[38] ), .D(\R_DATA_TEMPR27[38] ), .Y(
        OR4_341_Y));
    OR4 OR4_776 (.A(\R_DATA_TEMPR24[24] ), .B(\R_DATA_TEMPR25[24] ), 
        .C(\R_DATA_TEMPR26[24] ), .D(\R_DATA_TEMPR27[24] ), .Y(
        OR4_776_Y));
    OR4 OR4_763 (.A(\R_DATA_TEMPR36[2] ), .B(\R_DATA_TEMPR37[2] ), .C(
        \R_DATA_TEMPR38[2] ), .D(\R_DATA_TEMPR39[2] ), .Y(OR4_763_Y));
    OR4 OR4_264 (.A(OR4_571_Y), .B(OR4_40_Y), .C(OR4_384_Y), .D(
        OR4_713_Y), .Y(OR4_264_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%7%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R7C0 (.A_DOUT({
        \R_DATA_TEMPR7[39] , \R_DATA_TEMPR7[38] , \R_DATA_TEMPR7[37] , 
        \R_DATA_TEMPR7[36] , \R_DATA_TEMPR7[35] , \R_DATA_TEMPR7[34] , 
        \R_DATA_TEMPR7[33] , \R_DATA_TEMPR7[32] , \R_DATA_TEMPR7[31] , 
        \R_DATA_TEMPR7[30] , \R_DATA_TEMPR7[29] , \R_DATA_TEMPR7[28] , 
        \R_DATA_TEMPR7[27] , \R_DATA_TEMPR7[26] , \R_DATA_TEMPR7[25] , 
        \R_DATA_TEMPR7[24] , \R_DATA_TEMPR7[23] , \R_DATA_TEMPR7[22] , 
        \R_DATA_TEMPR7[21] , \R_DATA_TEMPR7[20] }), .B_DOUT({
        \R_DATA_TEMPR7[19] , \R_DATA_TEMPR7[18] , \R_DATA_TEMPR7[17] , 
        \R_DATA_TEMPR7[16] , \R_DATA_TEMPR7[15] , \R_DATA_TEMPR7[14] , 
        \R_DATA_TEMPR7[13] , \R_DATA_TEMPR7[12] , \R_DATA_TEMPR7[11] , 
        \R_DATA_TEMPR7[10] , \R_DATA_TEMPR7[9] , \R_DATA_TEMPR7[8] , 
        \R_DATA_TEMPR7[7] , \R_DATA_TEMPR7[6] , \R_DATA_TEMPR7[5] , 
        \R_DATA_TEMPR7[4] , \R_DATA_TEMPR7[3] , \R_DATA_TEMPR7[2] , 
        \R_DATA_TEMPR7[1] , \R_DATA_TEMPR7[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[7][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_656 (.A(OR4_237_Y), .B(OR4_258_Y), .C(OR4_243_Y), .D(
        OR4_622_Y), .Y(OR4_656_Y));
    OR4 OR4_440 (.A(\R_DATA_TEMPR28[12] ), .B(\R_DATA_TEMPR29[12] ), 
        .C(\R_DATA_TEMPR30[12] ), .D(\R_DATA_TEMPR31[12] ), .Y(
        OR4_440_Y));
    OR4 OR4_293 (.A(\R_DATA_TEMPR20[35] ), .B(\R_DATA_TEMPR21[35] ), 
        .C(\R_DATA_TEMPR22[35] ), .D(\R_DATA_TEMPR23[35] ), .Y(
        OR4_293_Y));
    OR4 OR4_388 (.A(\R_DATA_TEMPR28[37] ), .B(\R_DATA_TEMPR29[37] ), 
        .C(\R_DATA_TEMPR30[37] ), .D(\R_DATA_TEMPR31[37] ), .Y(
        OR4_388_Y));
    OR4 OR4_115 (.A(\R_DATA_TEMPR36[21] ), .B(\R_DATA_TEMPR37[21] ), 
        .C(\R_DATA_TEMPR38[21] ), .D(\R_DATA_TEMPR39[21] ), .Y(
        OR4_115_Y));
    OR4 OR4_66 (.A(\R_DATA_TEMPR48[23] ), .B(\R_DATA_TEMPR49[23] ), .C(
        \R_DATA_TEMPR50[23] ), .D(\R_DATA_TEMPR51[23] ), .Y(OR4_66_Y));
    OR4 OR4_417 (.A(OR4_629_Y), .B(OR4_504_Y), .C(OR4_776_Y), .D(
        OR4_476_Y), .Y(OR4_417_Y));
    OR4 OR4_433 (.A(\R_DATA_TEMPR44[17] ), .B(\R_DATA_TEMPR45[17] ), 
        .C(\R_DATA_TEMPR46[17] ), .D(\R_DATA_TEMPR47[17] ), .Y(
        OR4_433_Y));
    OR4 OR4_631 (.A(\R_DATA_TEMPR40[32] ), .B(\R_DATA_TEMPR41[32] ), 
        .C(\R_DATA_TEMPR42[32] ), .D(\R_DATA_TEMPR43[32] ), .Y(
        OR4_631_Y));
    OR4 OR4_365 (.A(\R_DATA_TEMPR0[5] ), .B(\R_DATA_TEMPR1[5] ), .C(
        \R_DATA_TEMPR2[5] ), .D(\R_DATA_TEMPR3[5] ), .Y(OR4_365_Y));
    OR4 OR4_238 (.A(\R_DATA_TEMPR56[17] ), .B(\R_DATA_TEMPR57[17] ), 
        .C(\R_DATA_TEMPR58[17] ), .D(\R_DATA_TEMPR59[17] ), .Y(
        OR4_238_Y));
    OR4 OR4_189 (.A(OR4_508_Y), .B(OR4_784_Y), .C(OR4_322_Y), .D(
        OR4_650_Y), .Y(OR4_189_Y));
    OR4 OR4_0 (.A(OR4_283_Y), .B(OR4_410_Y), .C(OR4_408_Y), .D(
        OR4_541_Y), .Y(OR4_0_Y));
    OR4 OR4_207 (.A(\R_DATA_TEMPR20[6] ), .B(\R_DATA_TEMPR21[6] ), .C(
        \R_DATA_TEMPR22[6] ), .D(\R_DATA_TEMPR23[6] ), .Y(OR4_207_Y));
    OR4 OR4_215 (.A(\R_DATA_TEMPR0[15] ), .B(\R_DATA_TEMPR1[15] ), .C(
        \R_DATA_TEMPR2[15] ), .D(\R_DATA_TEMPR3[15] ), .Y(OR4_215_Y));
    OR4 OR4_107 (.A(\R_DATA_TEMPR44[10] ), .B(\R_DATA_TEMPR45[10] ), 
        .C(\R_DATA_TEMPR46[10] ), .D(\R_DATA_TEMPR47[10] ), .Y(
        OR4_107_Y));
    OR4 OR4_277 (.A(\R_DATA_TEMPR12[3] ), .B(\R_DATA_TEMPR13[3] ), .C(
        \R_DATA_TEMPR14[3] ), .D(\R_DATA_TEMPR15[3] ), .Y(OR4_277_Y));
    OR4 OR4_698 (.A(\R_DATA_TEMPR52[15] ), .B(\R_DATA_TEMPR53[15] ), 
        .C(\R_DATA_TEMPR54[15] ), .D(\R_DATA_TEMPR55[15] ), .Y(
        OR4_698_Y));
    OR4 OR4_95 (.A(\R_DATA_TEMPR56[4] ), .B(\R_DATA_TEMPR57[4] ), .C(
        \R_DATA_TEMPR58[4] ), .D(\R_DATA_TEMPR59[4] ), .Y(OR4_95_Y));
    OR4 OR4_177 (.A(\R_DATA_TEMPR36[1] ), .B(\R_DATA_TEMPR37[1] ), .C(
        \R_DATA_TEMPR38[1] ), .D(\R_DATA_TEMPR39[1] ), .Y(OR4_177_Y));
    OR4 \OR4_R_DATA[34]  (.A(OR4_141_Y), .B(OR4_667_Y), .C(OR4_268_Y), 
        .D(OR4_603_Y), .Y(R_DATA[34]));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[14]  (.A(CFG3_1_Y), .B(CFG2_1_Y)
        , .Y(\BLKY2[14] ));
    OR4 OR4_762 (.A(OR4_102_Y), .B(OR4_576_Y), .C(OR4_737_Y), .D(
        OR4_343_Y), .Y(OR4_762_Y));
    OR4 OR4_349 (.A(\R_DATA_TEMPR28[1] ), .B(\R_DATA_TEMPR29[1] ), .C(
        \R_DATA_TEMPR30[1] ), .D(\R_DATA_TEMPR31[1] ), .Y(OR4_349_Y));
    OR4 OR4_692 (.A(OR4_561_Y), .B(OR4_730_Y), .C(OR4_19_Y), .D(
        OR4_607_Y), .Y(OR4_692_Y));
    OR4 OR4_703 (.A(\R_DATA_TEMPR8[3] ), .B(\R_DATA_TEMPR9[3] ), .C(
        \R_DATA_TEMPR10[3] ), .D(\R_DATA_TEMPR11[3] ), .Y(OR4_703_Y));
    OR4 OR4_223 (.A(\R_DATA_TEMPR40[37] ), .B(\R_DATA_TEMPR41[37] ), 
        .C(\R_DATA_TEMPR42[37] ), .D(\R_DATA_TEMPR43[37] ), .Y(
        OR4_223_Y));
    OR4 OR4_204 (.A(\R_DATA_TEMPR44[35] ), .B(\R_DATA_TEMPR45[35] ), 
        .C(\R_DATA_TEMPR46[35] ), .D(\R_DATA_TEMPR47[35] ), .Y(
        OR4_204_Y));
    OR4 OR4_354 (.A(OR4_366_Y), .B(OR4_520_Y), .C(OR4_254_Y), .D(
        OR4_670_Y), .Y(OR4_354_Y));
    OR4 OR4_773 (.A(\R_DATA_TEMPR28[29] ), .B(\R_DATA_TEMPR29[29] ), 
        .C(\R_DATA_TEMPR30[29] ), .D(\R_DATA_TEMPR31[29] ), .Y(
        OR4_773_Y));
    OR4 OR4_665 (.A(\R_DATA_TEMPR20[16] ), .B(\R_DATA_TEMPR21[16] ), 
        .C(\R_DATA_TEMPR22[16] ), .D(\R_DATA_TEMPR23[16] ), .Y(
        OR4_665_Y));
    OR4 OR4_413 (.A(OR4_271_Y), .B(OR4_382_Y), .C(OR4_474_Y), .D(
        OR4_434_Y), .Y(OR4_413_Y));
    OR4 OR4_611 (.A(\R_DATA_TEMPR4[25] ), .B(\R_DATA_TEMPR5[25] ), .C(
        \R_DATA_TEMPR6[25] ), .D(\R_DATA_TEMPR7[25] ), .Y(OR4_611_Y));
    OR4 OR4_151 (.A(\R_DATA_TEMPR8[28] ), .B(\R_DATA_TEMPR9[28] ), .C(
        \R_DATA_TEMPR10[28] ), .D(\R_DATA_TEMPR11[28] ), .Y(OR4_151_Y));
    OR4 OR4_274 (.A(\R_DATA_TEMPR24[29] ), .B(\R_DATA_TEMPR25[29] ), 
        .C(\R_DATA_TEMPR26[29] ), .D(\R_DATA_TEMPR27[29] ), .Y(
        OR4_274_Y));
    OR4 OR4_218 (.A(OR4_236_Y), .B(OR4_793_Y), .C(OR4_10_Y), .D(
        OR4_137_Y), .Y(OR4_218_Y));
    OR4 \OR4_R_DATA[22]  (.A(OR4_512_Y), .B(OR4_485_Y), .C(OR4_377_Y), 
        .D(OR4_18_Y), .Y(R_DATA[22]));
    OR4 OR4_60 (.A(OR4_315_Y), .B(OR4_63_Y), .C(OR4_98_Y), .D(
        OR4_468_Y), .Y(OR4_60_Y));
    OR4 OR4_531 (.A(\R_DATA_TEMPR8[2] ), .B(\R_DATA_TEMPR9[2] ), .C(
        \R_DATA_TEMPR10[2] ), .D(\R_DATA_TEMPR11[2] ), .Y(OR4_531_Y));
    OR4 OR4_67 (.A(\R_DATA_TEMPR40[26] ), .B(\R_DATA_TEMPR41[26] ), .C(
        \R_DATA_TEMPR42[26] ), .D(\R_DATA_TEMPR43[26] ), .Y(OR4_67_Y));
    OR4 OR4_785 (.A(OR4_84_Y), .B(OR4_246_Y), .C(OR4_360_Y), .D(
        OR4_275_Y), .Y(OR4_785_Y));
    OR4 OR4_687 (.A(\R_DATA_TEMPR0[23] ), .B(\R_DATA_TEMPR1[23] ), .C(
        \R_DATA_TEMPR2[23] ), .D(\R_DATA_TEMPR3[23] ), .Y(OR4_687_Y));
    OR4 OR4_305 (.A(\R_DATA_TEMPR60[27] ), .B(\R_DATA_TEMPR61[27] ), 
        .C(\R_DATA_TEMPR62[27] ), .D(\R_DATA_TEMPR63[27] ), .Y(
        OR4_305_Y));
    OR4 OR4_451 (.A(\R_DATA_TEMPR4[26] ), .B(\R_DATA_TEMPR5[26] ), .C(
        \R_DATA_TEMPR6[26] ), .D(\R_DATA_TEMPR7[26] ), .Y(OR4_451_Y));
    OR4 OR4_786 (.A(\R_DATA_TEMPR4[33] ), .B(\R_DATA_TEMPR5[33] ), .C(
        \R_DATA_TEMPR6[33] ), .D(\R_DATA_TEMPR7[33] ), .Y(OR4_786_Y));
    OR4 OR4_458 (.A(\R_DATA_TEMPR20[17] ), .B(\R_DATA_TEMPR21[17] ), 
        .C(\R_DATA_TEMPR22[17] ), .D(\R_DATA_TEMPR23[17] ), .Y(
        OR4_458_Y));
    OR4 OR4_628 (.A(\R_DATA_TEMPR4[0] ), .B(\R_DATA_TEMPR5[0] ), .C(
        \R_DATA_TEMPR6[0] ), .D(\R_DATA_TEMPR7[0] ), .Y(OR4_628_Y));
    OR4 OR4_375 (.A(OR4_438_Y), .B(OR4_197_Y), .C(OR4_221_Y), .D(
        OR4_395_Y), .Y(OR4_375_Y));
    OR4 OR4_749 (.A(OR4_113_Y), .B(OR4_680_Y), .C(OR4_133_Y), .D(
        OR4_364_Y), .Y(OR4_749_Y));
    OR4 OR4_660 (.A(OR4_636_Y), .B(OR4_628_Y), .C(OR4_572_Y), .D(
        OR4_781_Y), .Y(OR4_660_Y));
    OR4 OR4_622 (.A(\R_DATA_TEMPR28[18] ), .B(\R_DATA_TEMPR29[18] ), 
        .C(\R_DATA_TEMPR30[18] ), .D(\R_DATA_TEMPR31[18] ), .Y(
        OR4_622_Y));
    OR4 OR4_232 (.A(\R_DATA_TEMPR4[39] ), .B(\R_DATA_TEMPR5[39] ), .C(
        \R_DATA_TEMPR6[39] ), .D(\R_DATA_TEMPR7[39] ), .Y(OR4_232_Y));
    CFG3 #( .INIT(8'h20) )  CFG3_6 (.A(R_ADDR[13]), .B(R_ADDR[12]), .C(
        R_ADDR[11]), .Y(CFG3_6_Y));
    OR4 \OR4_R_DATA[15]  (.A(OR4_697_Y), .B(OR4_287_Y), .C(OR4_586_Y), 
        .D(OR4_363_Y), .Y(R_DATA[15]));
    OR4 OR4_543 (.A(\R_DATA_TEMPR56[35] ), .B(\R_DATA_TEMPR57[35] ), 
        .C(\R_DATA_TEMPR58[35] ), .D(\R_DATA_TEMPR59[35] ), .Y(
        OR4_543_Y));
    OR4 OR4_45 (.A(\R_DATA_TEMPR32[14] ), .B(\R_DATA_TEMPR33[14] ), .C(
        \R_DATA_TEMPR34[14] ), .D(\R_DATA_TEMPR35[14] ), .Y(OR4_45_Y));
    OR4 OR4_367 (.A(\R_DATA_TEMPR60[19] ), .B(\R_DATA_TEMPR61[19] ), 
        .C(\R_DATA_TEMPR62[19] ), .D(\R_DATA_TEMPR63[19] ), .Y(
        OR4_367_Y));
    OR4 OR4_160 (.A(\R_DATA_TEMPR12[8] ), .B(\R_DATA_TEMPR13[8] ), .C(
        \R_DATA_TEMPR14[8] ), .D(\R_DATA_TEMPR15[8] ), .Y(OR4_160_Y));
    OR4 OR4_702 (.A(\R_DATA_TEMPR4[9] ), .B(\R_DATA_TEMPR5[9] ), .C(
        \R_DATA_TEMPR6[9] ), .D(\R_DATA_TEMPR7[9] ), .Y(OR4_702_Y));
    OR4 OR4_559 (.A(\R_DATA_TEMPR8[12] ), .B(\R_DATA_TEMPR9[12] ), .C(
        \R_DATA_TEMPR10[12] ), .D(\R_DATA_TEMPR11[12] ), .Y(OR4_559_Y));
    OR4 OR4_550 (.A(\R_DATA_TEMPR56[13] ), .B(\R_DATA_TEMPR57[13] ), 
        .C(\R_DATA_TEMPR58[13] ), .D(\R_DATA_TEMPR59[13] ), .Y(
        OR4_550_Y));
    OR4 \OR4_R_DATA[23]  (.A(OR4_425_Y), .B(OR4_217_Y), .C(OR4_179_Y), 
        .D(OR4_155_Y), .Y(R_DATA[23]));
    OR4 OR4_330 (.A(\R_DATA_TEMPR4[22] ), .B(\R_DATA_TEMPR5[22] ), .C(
        \R_DATA_TEMPR6[22] ), .D(\R_DATA_TEMPR7[22] ), .Y(OR4_330_Y));
    OR4 OR4_772 (.A(\R_DATA_TEMPR0[7] ), .B(\R_DATA_TEMPR1[7] ), .C(
        \R_DATA_TEMPR2[7] ), .D(\R_DATA_TEMPR3[7] ), .Y(OR4_772_Y));
    OR4 OR4_768 (.A(OR4_555_Y), .B(OR4_432_Y), .C(OR4_297_Y), .D(
        OR4_305_Y), .Y(OR4_768_Y));
    OR4 OR4_605 (.A(\R_DATA_TEMPR56[34] ), .B(\R_DATA_TEMPR57[34] ), 
        .C(\R_DATA_TEMPR58[34] ), .D(\R_DATA_TEMPR59[34] ), .Y(
        OR4_605_Y));
    OR4 OR4_511 (.A(\R_DATA_TEMPR36[6] ), .B(\R_DATA_TEMPR37[6] ), .C(
        \R_DATA_TEMPR38[6] ), .D(\R_DATA_TEMPR39[6] ), .Y(OR4_511_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%14%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R14C0 (
        .A_DOUT({\R_DATA_TEMPR14[39] , \R_DATA_TEMPR14[38] , 
        \R_DATA_TEMPR14[37] , \R_DATA_TEMPR14[36] , 
        \R_DATA_TEMPR14[35] , \R_DATA_TEMPR14[34] , 
        \R_DATA_TEMPR14[33] , \R_DATA_TEMPR14[32] , 
        \R_DATA_TEMPR14[31] , \R_DATA_TEMPR14[30] , 
        \R_DATA_TEMPR14[29] , \R_DATA_TEMPR14[28] , 
        \R_DATA_TEMPR14[27] , \R_DATA_TEMPR14[26] , 
        \R_DATA_TEMPR14[25] , \R_DATA_TEMPR14[24] , 
        \R_DATA_TEMPR14[23] , \R_DATA_TEMPR14[22] , 
        \R_DATA_TEMPR14[21] , \R_DATA_TEMPR14[20] }), .B_DOUT({
        \R_DATA_TEMPR14[19] , \R_DATA_TEMPR14[18] , 
        \R_DATA_TEMPR14[17] , \R_DATA_TEMPR14[16] , 
        \R_DATA_TEMPR14[15] , \R_DATA_TEMPR14[14] , 
        \R_DATA_TEMPR14[13] , \R_DATA_TEMPR14[12] , 
        \R_DATA_TEMPR14[11] , \R_DATA_TEMPR14[10] , 
        \R_DATA_TEMPR14[9] , \R_DATA_TEMPR14[8] , \R_DATA_TEMPR14[7] , 
        \R_DATA_TEMPR14[6] , \R_DATA_TEMPR14[5] , \R_DATA_TEMPR14[4] , 
        \R_DATA_TEMPR14[3] , \R_DATA_TEMPR14[2] , \R_DATA_TEMPR14[1] , 
        \R_DATA_TEMPR14[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_696 (.A(OR4_126_Y), .B(OR4_547_Y), .C(OR4_13_Y), .D(
        OR4_521_Y), .Y(OR4_696_Y));
    OR4 OR4_675 (.A(OR4_131_Y), .B(OR4_786_Y), .C(OR4_769_Y), .D(
        OR4_453_Y), .Y(OR4_675_Y));
    OR4 OR4_287 (.A(OR4_771_Y), .B(OR4_184_Y), .C(OR4_173_Y), .D(
        OR4_553_Y), .Y(OR4_287_Y));
    OR4 OR4_86 (.A(\R_DATA_TEMPR12[36] ), .B(\R_DATA_TEMPR13[36] ), .C(
        \R_DATA_TEMPR14[36] ), .D(\R_DATA_TEMPR15[36] ), .Y(OR4_86_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[4]  (.A(CFG3_3_Y), .B(CFG2_2_Y), 
        .Y(\BLKX2[4] ));
    OR4 OR4_33 (.A(OR4_153_Y), .B(OR4_139_Y), .C(OR4_124_Y), .D(
        OR4_514_Y), .Y(OR4_33_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[10]  (.A(CFG3_0_Y), .B(CFG2_1_Y)
        , .Y(\BLKY2[10] ));
    OR4 OR4_168 (.A(\R_DATA_TEMPR0[27] ), .B(\R_DATA_TEMPR1[27] ), .C(
        \R_DATA_TEMPR2[27] ), .D(\R_DATA_TEMPR3[27] ), .Y(OR4_168_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%1%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R1C0 (.A_DOUT({
        \R_DATA_TEMPR1[39] , \R_DATA_TEMPR1[38] , \R_DATA_TEMPR1[37] , 
        \R_DATA_TEMPR1[36] , \R_DATA_TEMPR1[35] , \R_DATA_TEMPR1[34] , 
        \R_DATA_TEMPR1[33] , \R_DATA_TEMPR1[32] , \R_DATA_TEMPR1[31] , 
        \R_DATA_TEMPR1[30] , \R_DATA_TEMPR1[29] , \R_DATA_TEMPR1[28] , 
        \R_DATA_TEMPR1[27] , \R_DATA_TEMPR1[26] , \R_DATA_TEMPR1[25] , 
        \R_DATA_TEMPR1[24] , \R_DATA_TEMPR1[23] , \R_DATA_TEMPR1[22] , 
        \R_DATA_TEMPR1[21] , \R_DATA_TEMPR1[20] }), .B_DOUT({
        \R_DATA_TEMPR1[19] , \R_DATA_TEMPR1[18] , \R_DATA_TEMPR1[17] , 
        \R_DATA_TEMPR1[16] , \R_DATA_TEMPR1[15] , \R_DATA_TEMPR1[14] , 
        \R_DATA_TEMPR1[13] , \R_DATA_TEMPR1[12] , \R_DATA_TEMPR1[11] , 
        \R_DATA_TEMPR1[10] , \R_DATA_TEMPR1[9] , \R_DATA_TEMPR1[8] , 
        \R_DATA_TEMPR1[7] , \R_DATA_TEMPR1[6] , \R_DATA_TEMPR1[5] , 
        \R_DATA_TEMPR1[4] , \R_DATA_TEMPR1[3] , \R_DATA_TEMPR1[2] , 
        \R_DATA_TEMPR1[1] , \R_DATA_TEMPR1[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[1][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_187 (.A(OR4_103_Y), .B(OR4_369_Y), .C(OR4_195_Y), .D(
        OR4_192_Y), .Y(OR4_187_Y));
    OR4 OR4_212 (.A(\R_DATA_TEMPR20[3] ), .B(\R_DATA_TEMPR21[3] ), .C(
        \R_DATA_TEMPR22[3] ), .D(\R_DATA_TEMPR23[3] ), .Y(OR4_212_Y));
    OR4 OR4_353 (.A(\R_DATA_TEMPR20[38] ), .B(\R_DATA_TEMPR21[38] ), 
        .C(\R_DATA_TEMPR22[38] ), .D(\R_DATA_TEMPR23[38] ), .Y(
        OR4_353_Y));
    OR4 OR4_750 (.A(\R_DATA_TEMPR40[29] ), .B(\R_DATA_TEMPR41[29] ), 
        .C(\R_DATA_TEMPR42[29] ), .D(\R_DATA_TEMPR43[29] ), .Y(
        OR4_750_Y));
    OR4 OR4_783 (.A(\R_DATA_TEMPR0[30] ), .B(\R_DATA_TEMPR1[30] ), .C(
        \R_DATA_TEMPR2[30] ), .D(\R_DATA_TEMPR3[30] ), .Y(OR4_783_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[2]  (.A(CFG3_0_Y), .B(CFG2_0_Y), 
        .Y(\BLKY2[2] ));
    OR4 OR4_600 (.A(\R_DATA_TEMPR8[10] ), .B(\R_DATA_TEMPR9[10] ), .C(
        \R_DATA_TEMPR10[10] ), .D(\R_DATA_TEMPR11[10] ), .Y(OR4_600_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%11%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R11C0 (
        .A_DOUT({\R_DATA_TEMPR11[39] , \R_DATA_TEMPR11[38] , 
        \R_DATA_TEMPR11[37] , \R_DATA_TEMPR11[36] , 
        \R_DATA_TEMPR11[35] , \R_DATA_TEMPR11[34] , 
        \R_DATA_TEMPR11[33] , \R_DATA_TEMPR11[32] , 
        \R_DATA_TEMPR11[31] , \R_DATA_TEMPR11[30] , 
        \R_DATA_TEMPR11[29] , \R_DATA_TEMPR11[28] , 
        \R_DATA_TEMPR11[27] , \R_DATA_TEMPR11[26] , 
        \R_DATA_TEMPR11[25] , \R_DATA_TEMPR11[24] , 
        \R_DATA_TEMPR11[23] , \R_DATA_TEMPR11[22] , 
        \R_DATA_TEMPR11[21] , \R_DATA_TEMPR11[20] }), .B_DOUT({
        \R_DATA_TEMPR11[19] , \R_DATA_TEMPR11[18] , 
        \R_DATA_TEMPR11[17] , \R_DATA_TEMPR11[16] , 
        \R_DATA_TEMPR11[15] , \R_DATA_TEMPR11[14] , 
        \R_DATA_TEMPR11[13] , \R_DATA_TEMPR11[12] , 
        \R_DATA_TEMPR11[11] , \R_DATA_TEMPR11[10] , 
        \R_DATA_TEMPR11[9] , \R_DATA_TEMPR11[8] , \R_DATA_TEMPR11[7] , 
        \R_DATA_TEMPR11[6] , \R_DATA_TEMPR11[5] , \R_DATA_TEMPR11[4] , 
        \R_DATA_TEMPR11[3] , \R_DATA_TEMPR11[2] , \R_DATA_TEMPR11[1] , 
        \R_DATA_TEMPR11[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[2] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_452 (.A(\R_DATA_TEMPR36[5] ), .B(\R_DATA_TEMPR37[5] ), .C(
        \R_DATA_TEMPR38[5] ), .D(\R_DATA_TEMPR39[5] ), .Y(OR4_452_Y));
    OR4 OR4_284 (.A(\R_DATA_TEMPR24[35] ), .B(\R_DATA_TEMPR25[35] ), 
        .C(\R_DATA_TEMPR26[35] ), .D(\R_DATA_TEMPR27[35] ), .Y(
        OR4_284_Y));
    OR4 OR4_310 (.A(OR4_691_Y), .B(OR4_451_Y), .C(OR4_495_Y), .D(
        OR4_643_Y), .Y(OR4_310_Y));
    OR4 OR4_5 (.A(OR4_596_Y), .B(OR4_71_Y), .C(OR4_463_Y), .D(
        OR4_589_Y), .Y(OR4_5_Y));
    OR4 OR4_670 (.A(\R_DATA_TEMPR44[3] ), .B(\R_DATA_TEMPR45[3] ), .C(
        \R_DATA_TEMPR46[3] ), .D(\R_DATA_TEMPR47[3] ), .Y(OR4_670_Y));
    OR4 OR4_459 (.A(OR4_387_Y), .B(OR4_272_Y), .C(OR4_116_Y), .D(
        OR4_506_Y), .Y(OR4_459_Y));
    OR4 OR4_307 (.A(\R_DATA_TEMPR40[39] ), .B(\R_DATA_TEMPR41[39] ), 
        .C(\R_DATA_TEMPR42[39] ), .D(\R_DATA_TEMPR43[39] ), .Y(
        OR4_307_Y));
    OR4 OR4_100 (.A(OR4_168_Y), .B(OR4_615_Y), .C(OR4_110_Y), .D(
        OR4_499_Y), .Y(OR4_100_Y));
    OR4 OR4_99 (.A(\R_DATA_TEMPR28[8] ), .B(\R_DATA_TEMPR29[8] ), .C(
        \R_DATA_TEMPR30[8] ), .D(\R_DATA_TEMPR31[8] ), .Y(OR4_99_Y));
    OR4 OR4_156 (.A(\R_DATA_TEMPR44[15] ), .B(\R_DATA_TEMPR45[15] ), 
        .C(\R_DATA_TEMPR46[15] ), .D(\R_DATA_TEMPR47[15] ), .Y(
        OR4_156_Y));
    OR4 OR4_535 (.A(\R_DATA_TEMPR24[19] ), .B(\R_DATA_TEMPR25[19] ), 
        .C(\R_DATA_TEMPR26[19] ), .D(\R_DATA_TEMPR27[19] ), .Y(
        OR4_535_Y));
    OR4 OR4_68 (.A(\R_DATA_TEMPR16[34] ), .B(\R_DATA_TEMPR17[34] ), .C(
        \R_DATA_TEMPR18[34] ), .D(\R_DATA_TEMPR19[34] ), .Y(OR4_68_Y));
    OR4 OR4_377 (.A(OR4_416_Y), .B(OR4_695_Y), .C(OR4_289_Y), .D(
        OR4_409_Y), .Y(OR4_377_Y));
    OR4 OR4_170 (.A(OR4_240_Y), .B(OR4_678_Y), .C(OR4_185_Y), .D(
        OR4_562_Y), .Y(OR4_170_Y));
    OR4 OR4_708 (.A(\R_DATA_TEMPR24[25] ), .B(\R_DATA_TEMPR25[25] ), 
        .C(\R_DATA_TEMPR26[25] ), .D(\R_DATA_TEMPR27[25] ), .Y(
        OR4_708_Y));
    OR4 OR4_626 (.A(\R_DATA_TEMPR60[29] ), .B(\R_DATA_TEMPR61[29] ), 
        .C(\R_DATA_TEMPR62[29] ), .D(\R_DATA_TEMPR63[29] ), .Y(
        OR4_626_Y));
    OR4 OR4_31 (.A(OR4_260_Y), .B(OR4_172_Y), .C(OR4_238_Y), .D(
        OR4_42_Y), .Y(OR4_31_Y));
    OR4 OR4_633 (.A(OR4_142_Y), .B(OR4_611_Y), .C(OR4_646_Y), .D(
        OR4_256_Y), .Y(OR4_633_Y));
    OR4 \OR4_R_DATA[31]  (.A(OR4_188_Y), .B(OR4_146_Y), .C(OR4_159_Y), 
        .D(OR4_712_Y), .Y(R_DATA[31]));
    OR4 OR4_385 (.A(\R_DATA_TEMPR24[9] ), .B(\R_DATA_TEMPR25[9] ), .C(
        \R_DATA_TEMPR26[9] ), .D(\R_DATA_TEMPR27[9] ), .Y(OR4_385_Y));
    OR4 OR4_778 (.A(OR4_329_Y), .B(OR4_248_Y), .C(OR4_739_Y), .D(
        OR4_204_Y), .Y(OR4_778_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[15]  (.A(CFG3_15_Y), .B(
        CFG2_3_Y), .Y(\BLKX2[15] ));
    OR4 OR4_243 (.A(\R_DATA_TEMPR24[18] ), .B(\R_DATA_TEMPR25[18] ), 
        .C(\R_DATA_TEMPR26[18] ), .D(\R_DATA_TEMPR27[18] ), .Y(
        OR4_243_Y));
    OR4 OR4_394 (.A(\R_DATA_TEMPR4[12] ), .B(\R_DATA_TEMPR5[12] ), .C(
        \R_DATA_TEMPR6[12] ), .D(\R_DATA_TEMPR7[12] ), .Y(OR4_394_Y));
    OR4 OR4_358 (.A(\R_DATA_TEMPR4[20] ), .B(\R_DATA_TEMPR5[20] ), .C(
        \R_DATA_TEMPR6[20] ), .D(\R_DATA_TEMPR7[20] ), .Y(OR4_358_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%20%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R20C0 (
        .A_DOUT({\R_DATA_TEMPR20[39] , \R_DATA_TEMPR20[38] , 
        \R_DATA_TEMPR20[37] , \R_DATA_TEMPR20[36] , 
        \R_DATA_TEMPR20[35] , \R_DATA_TEMPR20[34] , 
        \R_DATA_TEMPR20[33] , \R_DATA_TEMPR20[32] , 
        \R_DATA_TEMPR20[31] , \R_DATA_TEMPR20[30] , 
        \R_DATA_TEMPR20[29] , \R_DATA_TEMPR20[28] , 
        \R_DATA_TEMPR20[27] , \R_DATA_TEMPR20[26] , 
        \R_DATA_TEMPR20[25] , \R_DATA_TEMPR20[24] , 
        \R_DATA_TEMPR20[23] , \R_DATA_TEMPR20[22] , 
        \R_DATA_TEMPR20[21] , \R_DATA_TEMPR20[20] }), .B_DOUT({
        \R_DATA_TEMPR20[19] , \R_DATA_TEMPR20[18] , 
        \R_DATA_TEMPR20[17] , \R_DATA_TEMPR20[16] , 
        \R_DATA_TEMPR20[15] , \R_DATA_TEMPR20[14] , 
        \R_DATA_TEMPR20[13] , \R_DATA_TEMPR20[12] , 
        \R_DATA_TEMPR20[11] , \R_DATA_TEMPR20[10] , 
        \R_DATA_TEMPR20[9] , \R_DATA_TEMPR20[8] , \R_DATA_TEMPR20[7] , 
        \R_DATA_TEMPR20[6] , \R_DATA_TEMPR20[5] , \R_DATA_TEMPR20[4] , 
        \R_DATA_TEMPR20[3] , \R_DATA_TEMPR20[2] , \R_DATA_TEMPR20[1] , 
        \R_DATA_TEMPR20[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[5] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_80 (.A(OR4_661_Y), .B(OR4_575_Y), .C(OR4_647_Y), .D(
        OR4_46_Y), .Y(OR4_80_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R47C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%47%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R47C0 (
        .A_DOUT({\R_DATA_TEMPR47[39] , \R_DATA_TEMPR47[38] , 
        \R_DATA_TEMPR47[37] , \R_DATA_TEMPR47[36] , 
        \R_DATA_TEMPR47[35] , \R_DATA_TEMPR47[34] , 
        \R_DATA_TEMPR47[33] , \R_DATA_TEMPR47[32] , 
        \R_DATA_TEMPR47[31] , \R_DATA_TEMPR47[30] , 
        \R_DATA_TEMPR47[29] , \R_DATA_TEMPR47[28] , 
        \R_DATA_TEMPR47[27] , \R_DATA_TEMPR47[26] , 
        \R_DATA_TEMPR47[25] , \R_DATA_TEMPR47[24] , 
        \R_DATA_TEMPR47[23] , \R_DATA_TEMPR47[22] , 
        \R_DATA_TEMPR47[21] , \R_DATA_TEMPR47[20] }), .B_DOUT({
        \R_DATA_TEMPR47[19] , \R_DATA_TEMPR47[18] , 
        \R_DATA_TEMPR47[17] , \R_DATA_TEMPR47[16] , 
        \R_DATA_TEMPR47[15] , \R_DATA_TEMPR47[14] , 
        \R_DATA_TEMPR47[13] , \R_DATA_TEMPR47[12] , 
        \R_DATA_TEMPR47[11] , \R_DATA_TEMPR47[10] , 
        \R_DATA_TEMPR47[9] , \R_DATA_TEMPR47[8] , \R_DATA_TEMPR47[7] , 
        \R_DATA_TEMPR47[6] , \R_DATA_TEMPR47[5] , \R_DATA_TEMPR47[4] , 
        \R_DATA_TEMPR47[3] , \R_DATA_TEMPR47[2] , \R_DATA_TEMPR47[1] , 
        \R_DATA_TEMPR47[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[47][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[11] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[11] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_108 (.A(\R_DATA_TEMPR4[7] ), .B(\R_DATA_TEMPR5[7] ), .C(
        \R_DATA_TEMPR6[7] ), .D(\R_DATA_TEMPR7[7] ), .Y(OR4_108_Y));
    OR4 OR4_191 (.A(OR4_454_Y), .B(OR4_376_Y), .C(OR4_439_Y), .D(
        OR4_302_Y), .Y(OR4_191_Y));
    OR4 OR4_1 (.A(\R_DATA_TEMPR52[4] ), .B(\R_DATA_TEMPR53[4] ), .C(
        \R_DATA_TEMPR54[4] ), .D(\R_DATA_TEMPR55[4] ), .Y(OR4_1_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%29%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R29C0 (
        .A_DOUT({\R_DATA_TEMPR29[39] , \R_DATA_TEMPR29[38] , 
        \R_DATA_TEMPR29[37] , \R_DATA_TEMPR29[36] , 
        \R_DATA_TEMPR29[35] , \R_DATA_TEMPR29[34] , 
        \R_DATA_TEMPR29[33] , \R_DATA_TEMPR29[32] , 
        \R_DATA_TEMPR29[31] , \R_DATA_TEMPR29[30] , 
        \R_DATA_TEMPR29[29] , \R_DATA_TEMPR29[28] , 
        \R_DATA_TEMPR29[27] , \R_DATA_TEMPR29[26] , 
        \R_DATA_TEMPR29[25] , \R_DATA_TEMPR29[24] , 
        \R_DATA_TEMPR29[23] , \R_DATA_TEMPR29[22] , 
        \R_DATA_TEMPR29[21] , \R_DATA_TEMPR29[20] }), .B_DOUT({
        \R_DATA_TEMPR29[19] , \R_DATA_TEMPR29[18] , 
        \R_DATA_TEMPR29[17] , \R_DATA_TEMPR29[16] , 
        \R_DATA_TEMPR29[15] , \R_DATA_TEMPR29[14] , 
        \R_DATA_TEMPR29[13] , \R_DATA_TEMPR29[12] , 
        \R_DATA_TEMPR29[11] , \R_DATA_TEMPR29[10] , 
        \R_DATA_TEMPR29[9] , \R_DATA_TEMPR29[8] , \R_DATA_TEMPR29[7] , 
        \R_DATA_TEMPR29[6] , \R_DATA_TEMPR29[5] , \R_DATA_TEMPR29[4] , 
        \R_DATA_TEMPR29[3] , \R_DATA_TEMPR29[2] , \R_DATA_TEMPR29[1] , 
        \R_DATA_TEMPR29[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[7] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_87 (.A(\R_DATA_TEMPR16[20] ), .B(\R_DATA_TEMPR17[20] ), .C(
        \R_DATA_TEMPR18[20] ), .D(\R_DATA_TEMPR19[20] ), .Y(OR4_87_Y));
    OR4 \OR4_R_DATA[30]  (.A(OR4_36_Y), .B(OR4_224_Y), .C(OR4_581_Y), 
        .D(OR4_285_Y), .Y(R_DATA[30]));
    OR4 OR4_178 (.A(\R_DATA_TEMPR24[27] ), .B(\R_DATA_TEMPR25[27] ), 
        .C(\R_DATA_TEMPR26[27] ), .D(\R_DATA_TEMPR27[27] ), .Y(
        OR4_178_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[0]  (.A(CFG3_7_Y), .B(CFG2_2_Y), 
        .Y(\BLKX2[0] ));
    OR4 OR4_782 (.A(\R_DATA_TEMPR56[20] ), .B(\R_DATA_TEMPR57[20] ), 
        .C(\R_DATA_TEMPR58[20] ), .D(\R_DATA_TEMPR59[20] ), .Y(
        OR4_782_Y));
    OR4 OR4_159 (.A(OR4_437_Y), .B(OR4_348_Y), .C(OR4_50_Y), .D(
        OR4_313_Y), .Y(OR4_159_Y));
    OR4 OR4_491 (.A(\R_DATA_TEMPR56[26] ), .B(\R_DATA_TEMPR57[26] ), 
        .C(\R_DATA_TEMPR58[26] ), .D(\R_DATA_TEMPR59[26] ), .Y(
        OR4_491_Y));
    OR4 OR4_165 (.A(\R_DATA_TEMPR16[28] ), .B(\R_DATA_TEMPR17[28] ), 
        .C(\R_DATA_TEMPR18[28] ), .D(\R_DATA_TEMPR19[28] ), .Y(
        OR4_165_Y));
    OR4 OR4_133 (.A(\R_DATA_TEMPR24[0] ), .B(\R_DATA_TEMPR25[0] ), .C(
        \R_DATA_TEMPR26[0] ), .D(\R_DATA_TEMPR27[0] ), .Y(OR4_133_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%26%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R26C0 (
        .A_DOUT({\R_DATA_TEMPR26[39] , \R_DATA_TEMPR26[38] , 
        \R_DATA_TEMPR26[37] , \R_DATA_TEMPR26[36] , 
        \R_DATA_TEMPR26[35] , \R_DATA_TEMPR26[34] , 
        \R_DATA_TEMPR26[33] , \R_DATA_TEMPR26[32] , 
        \R_DATA_TEMPR26[31] , \R_DATA_TEMPR26[30] , 
        \R_DATA_TEMPR26[29] , \R_DATA_TEMPR26[28] , 
        \R_DATA_TEMPR26[27] , \R_DATA_TEMPR26[26] , 
        \R_DATA_TEMPR26[25] , \R_DATA_TEMPR26[24] , 
        \R_DATA_TEMPR26[23] , \R_DATA_TEMPR26[22] , 
        \R_DATA_TEMPR26[21] , \R_DATA_TEMPR26[20] }), .B_DOUT({
        \R_DATA_TEMPR26[19] , \R_DATA_TEMPR26[18] , 
        \R_DATA_TEMPR26[17] , \R_DATA_TEMPR26[16] , 
        \R_DATA_TEMPR26[15] , \R_DATA_TEMPR26[14] , 
        \R_DATA_TEMPR26[13] , \R_DATA_TEMPR26[12] , 
        \R_DATA_TEMPR26[11] , \R_DATA_TEMPR26[10] , 
        \R_DATA_TEMPR26[9] , \R_DATA_TEMPR26[8] , \R_DATA_TEMPR26[7] , 
        \R_DATA_TEMPR26[6] , \R_DATA_TEMPR26[5] , \R_DATA_TEMPR26[4] , 
        \R_DATA_TEMPR26[3] , \R_DATA_TEMPR26[2] , \R_DATA_TEMPR26[1] , 
        \R_DATA_TEMPR26[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[6] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[6] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_515 (.A(\R_DATA_TEMPR52[29] ), .B(\R_DATA_TEMPR53[29] ), 
        .C(\R_DATA_TEMPR54[29] ), .D(\R_DATA_TEMPR55[29] ), .Y(
        OR4_515_Y));
    OR4 OR4_498 (.A(\R_DATA_TEMPR12[35] ), .B(\R_DATA_TEMPR13[35] ), 
        .C(\R_DATA_TEMPR14[35] ), .D(\R_DATA_TEMPR15[35] ), .Y(
        OR4_498_Y));
    OR4 OR4_92 (.A(\R_DATA_TEMPR0[4] ), .B(\R_DATA_TEMPR1[4] ), .C(
        \R_DATA_TEMPR2[4] ), .D(\R_DATA_TEMPR3[4] ), .Y(OR4_92_Y));
    OR4 \OR4_R_DATA[36]  (.A(OR4_556_Y), .B(OR4_193_Y), .C(OR4_332_Y), 
        .D(OR4_375_Y), .Y(R_DATA[36]));
    OR4 OR4_467 (.A(OR4_772_Y), .B(OR4_108_Y), .C(OR4_583_Y), .D(
        OR4_493_Y), .Y(OR4_467_Y));
    OR4 OR4_648 (.A(\R_DATA_TEMPR32[7] ), .B(\R_DATA_TEMPR33[7] ), .C(
        \R_DATA_TEMPR34[7] ), .D(\R_DATA_TEMPR35[7] ), .Y(OR4_648_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%8%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R8C0 (.A_DOUT({
        \R_DATA_TEMPR8[39] , \R_DATA_TEMPR8[38] , \R_DATA_TEMPR8[37] , 
        \R_DATA_TEMPR8[36] , \R_DATA_TEMPR8[35] , \R_DATA_TEMPR8[34] , 
        \R_DATA_TEMPR8[33] , \R_DATA_TEMPR8[32] , \R_DATA_TEMPR8[31] , 
        \R_DATA_TEMPR8[30] , \R_DATA_TEMPR8[29] , \R_DATA_TEMPR8[28] , 
        \R_DATA_TEMPR8[27] , \R_DATA_TEMPR8[26] , \R_DATA_TEMPR8[25] , 
        \R_DATA_TEMPR8[24] , \R_DATA_TEMPR8[23] , \R_DATA_TEMPR8[22] , 
        \R_DATA_TEMPR8[21] , \R_DATA_TEMPR8[20] }), .B_DOUT({
        \R_DATA_TEMPR8[19] , \R_DATA_TEMPR8[18] , \R_DATA_TEMPR8[17] , 
        \R_DATA_TEMPR8[16] , \R_DATA_TEMPR8[15] , \R_DATA_TEMPR8[14] , 
        \R_DATA_TEMPR8[13] , \R_DATA_TEMPR8[12] , \R_DATA_TEMPR8[11] , 
        \R_DATA_TEMPR8[10] , \R_DATA_TEMPR8[9] , \R_DATA_TEMPR8[8] , 
        \R_DATA_TEMPR8[7] , \R_DATA_TEMPR8[6] , \R_DATA_TEMPR8[5] , 
        \R_DATA_TEMPR8[4] , \R_DATA_TEMPR8[3] , \R_DATA_TEMPR8[2] , 
        \R_DATA_TEMPR8[1] , \R_DATA_TEMPR8[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[8][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_685 (.A(\R_DATA_TEMPR32[39] ), .B(\R_DATA_TEMPR33[39] ), 
        .C(\R_DATA_TEMPR34[39] ), .D(\R_DATA_TEMPR35[39] ), .Y(
        OR4_685_Y));
    OR4 OR4_613 (.A(\R_DATA_TEMPR28[9] ), .B(\R_DATA_TEMPR29[9] ), .C(
        \R_DATA_TEMPR30[9] ), .D(\R_DATA_TEMPR31[9] ), .Y(OR4_613_Y));
    OR4 OR4_642 (.A(\R_DATA_TEMPR32[21] ), .B(\R_DATA_TEMPR33[21] ), 
        .C(\R_DATA_TEMPR34[21] ), .D(\R_DATA_TEMPR35[21] ), .Y(
        OR4_642_Y));
    CFG2 #( .INIT(4'h2) )  CFG2_0 (.A(R_EN), .B(R_ADDR[14]), .Y(
        CFG2_0_Y));
    OR4 OR4_324 (.A(\R_DATA_TEMPR44[1] ), .B(\R_DATA_TEMPR45[1] ), .C(
        \R_DATA_TEMPR46[1] ), .D(\R_DATA_TEMPR47[1] ), .Y(OR4_324_Y));
    OR4 OR4_265 (.A(\R_DATA_TEMPR32[17] ), .B(\R_DATA_TEMPR33[17] ), 
        .C(\R_DATA_TEMPR34[17] ), .D(\R_DATA_TEMPR35[17] ), .Y(
        OR4_265_Y));
    OR4 OR4_49 (.A(\R_DATA_TEMPR24[12] ), .B(\R_DATA_TEMPR25[12] ), .C(
        \R_DATA_TEMPR26[12] ), .D(\R_DATA_TEMPR27[12] ), .Y(OR4_49_Y));
    OR4 OR4_599 (.A(OR4_465_Y), .B(OR4_593_Y), .C(OR4_684_Y), .D(
        OR4_510_Y), .Y(OR4_599_Y));
    OR4 OR4_590 (.A(\R_DATA_TEMPR8[31] ), .B(\R_DATA_TEMPR9[31] ), .C(
        \R_DATA_TEMPR10[31] ), .D(\R_DATA_TEMPR11[31] ), .Y(OR4_590_Y));
    OR4 OR4_121 (.A(\R_DATA_TEMPR16[5] ), .B(\R_DATA_TEMPR17[5] ), .C(
        \R_DATA_TEMPR18[5] ), .D(\R_DATA_TEMPR19[5] ), .Y(OR4_121_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[5]  (.A(CFG3_14_Y), .B(CFG2_2_Y)
        , .Y(\BLKX2[5] ));
    OR4 \OR4_R_DATA[18]  (.A(OR4_760_Y), .B(OR4_656_Y), .C(OR4_298_Y), 
        .D(OR4_401_Y), .Y(R_DATA[18]));
    OR4 OR4_680 (.A(\R_DATA_TEMPR20[0] ), .B(\R_DATA_TEMPR21[0] ), .C(
        \R_DATA_TEMPR22[0] ), .D(\R_DATA_TEMPR23[0] ), .Y(OR4_680_Y));
    OR4 OR4_113 (.A(\R_DATA_TEMPR16[0] ), .B(\R_DATA_TEMPR17[0] ), .C(
        \R_DATA_TEMPR18[0] ), .D(\R_DATA_TEMPR19[0] ), .Y(OR4_113_Y));
    OR4 OR4_132 (.A(\R_DATA_TEMPR28[2] ), .B(\R_DATA_TEMPR29[2] ), .C(
        \R_DATA_TEMPR30[2] ), .D(\R_DATA_TEMPR31[2] ), .Y(OR4_132_Y));
    OR4 OR4_7 (.A(\R_DATA_TEMPR40[34] ), .B(\R_DATA_TEMPR41[34] ), .C(
        \R_DATA_TEMPR42[34] ), .D(\R_DATA_TEMPR43[34] ), .Y(OR4_7_Y));
    OR4 OR4_421 (.A(\R_DATA_TEMPR20[8] ), .B(\R_DATA_TEMPR21[8] ), .C(
        \R_DATA_TEMPR22[8] ), .D(\R_DATA_TEMPR23[8] ), .Y(OR4_421_Y));
    OR4 OR4_463 (.A(\R_DATA_TEMPR40[24] ), .B(\R_DATA_TEMPR41[24] ), 
        .C(\R_DATA_TEMPR42[24] ), .D(\R_DATA_TEMPR43[24] ), .Y(
        OR4_463_Y));
    OR4 OR4_755 (.A(\R_DATA_TEMPR0[16] ), .B(\R_DATA_TEMPR1[16] ), .C(
        \R_DATA_TEMPR2[16] ), .D(\R_DATA_TEMPR3[16] ), .Y(OR4_755_Y));
    OR4 OR4_661 (.A(\R_DATA_TEMPR48[12] ), .B(\R_DATA_TEMPR49[12] ), 
        .C(\R_DATA_TEMPR50[12] ), .D(\R_DATA_TEMPR51[12] ), .Y(
        OR4_661_Y));
    OR4 OR4_657 (.A(\R_DATA_TEMPR52[10] ), .B(\R_DATA_TEMPR53[10] ), 
        .C(\R_DATA_TEMPR54[10] ), .D(\R_DATA_TEMPR55[10] ), .Y(
        OR4_657_Y));
    OR4 OR4_428 (.A(\R_DATA_TEMPR40[36] ), .B(\R_DATA_TEMPR41[36] ), 
        .C(\R_DATA_TEMPR42[36] ), .D(\R_DATA_TEMPR43[36] ), .Y(
        OR4_428_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R61C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%61%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R61C0 (
        .A_DOUT({\R_DATA_TEMPR61[39] , \R_DATA_TEMPR61[38] , 
        \R_DATA_TEMPR61[37] , \R_DATA_TEMPR61[36] , 
        \R_DATA_TEMPR61[35] , \R_DATA_TEMPR61[34] , 
        \R_DATA_TEMPR61[33] , \R_DATA_TEMPR61[32] , 
        \R_DATA_TEMPR61[31] , \R_DATA_TEMPR61[30] , 
        \R_DATA_TEMPR61[29] , \R_DATA_TEMPR61[28] , 
        \R_DATA_TEMPR61[27] , \R_DATA_TEMPR61[26] , 
        \R_DATA_TEMPR61[25] , \R_DATA_TEMPR61[24] , 
        \R_DATA_TEMPR61[23] , \R_DATA_TEMPR61[22] , 
        \R_DATA_TEMPR61[21] , \R_DATA_TEMPR61[20] }), .B_DOUT({
        \R_DATA_TEMPR61[19] , \R_DATA_TEMPR61[18] , 
        \R_DATA_TEMPR61[17] , \R_DATA_TEMPR61[16] , 
        \R_DATA_TEMPR61[15] , \R_DATA_TEMPR61[14] , 
        \R_DATA_TEMPR61[13] , \R_DATA_TEMPR61[12] , 
        \R_DATA_TEMPR61[11] , \R_DATA_TEMPR61[10] , 
        \R_DATA_TEMPR61[9] , \R_DATA_TEMPR61[8] , \R_DATA_TEMPR61[7] , 
        \R_DATA_TEMPR61[6] , \R_DATA_TEMPR61[5] , \R_DATA_TEMPR61[4] , 
        \R_DATA_TEMPR61[3] , \R_DATA_TEMPR61[2] , \R_DATA_TEMPR61[1] , 
        \R_DATA_TEMPR61[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[61][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[15] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[15] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_756 (.A(\R_DATA_TEMPR0[39] ), .B(\R_DATA_TEMPR1[39] ), .C(
        \R_DATA_TEMPR2[39] ), .D(\R_DATA_TEMPR3[39] ), .Y(OR4_756_Y));
    OR4 OR4_268 (.A(OR4_389_Y), .B(OR4_309_Y), .C(OR4_7_Y), .D(
        OR4_276_Y), .Y(OR4_268_Y));
    OR4 OR4_387 (.A(\R_DATA_TEMPR48[21] ), .B(\R_DATA_TEMPR49[21] ), 
        .C(\R_DATA_TEMPR50[21] ), .D(\R_DATA_TEMPR51[21] ), .Y(
        OR4_387_Y));
    OR4 OR4_180 (.A(\R_DATA_TEMPR28[34] ), .B(\R_DATA_TEMPR29[34] ), 
        .C(\R_DATA_TEMPR30[34] ), .D(\R_DATA_TEMPR31[34] ), .Y(
        OR4_180_Y));
    OR4 OR4_105 (.A(\R_DATA_TEMPR44[2] ), .B(\R_DATA_TEMPR45[2] ), .C(
        \R_DATA_TEMPR46[2] ), .D(\R_DATA_TEMPR47[2] ), .Y(OR4_105_Y));
    OR4 OR4_788 (.A(\R_DATA_TEMPR48[15] ), .B(\R_DATA_TEMPR49[15] ), 
        .C(\R_DATA_TEMPR50[15] ), .D(\R_DATA_TEMPR51[15] ), .Y(
        OR4_788_Y));
    OR4 OR4_407 (.A(OR4_548_Y), .B(OR4_312_Y), .C(OR4_333_Y), .D(
        OR4_673_Y), .Y(OR4_407_Y));
    CFG3 #( .INIT(8'h80) )  CFG3_15 (.A(W_ADDR[13]), .B(W_ADDR[12]), 
        .C(W_ADDR[11]), .Y(CFG3_15_Y));
    OR4 OR4_175 (.A(\R_DATA_TEMPR48[9] ), .B(\R_DATA_TEMPR49[9] ), .C(
        \R_DATA_TEMPR50[9] ), .D(\R_DATA_TEMPR51[9] ), .Y(OR4_175_Y));
    OR4 OR4_393 (.A(\R_DATA_TEMPR0[35] ), .B(\R_DATA_TEMPR1[35] ), .C(
        \R_DATA_TEMPR2[35] ), .D(\R_DATA_TEMPR3[35] ), .Y(OR4_393_Y));
    OR4 OR4_790 (.A(\R_DATA_TEMPR32[15] ), .B(\R_DATA_TEMPR33[15] ), 
        .C(\R_DATA_TEMPR34[15] ), .D(\R_DATA_TEMPR35[15] ), .Y(
        OR4_790_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R50C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%50%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R50C0 (
        .A_DOUT({\R_DATA_TEMPR50[39] , \R_DATA_TEMPR50[38] , 
        \R_DATA_TEMPR50[37] , \R_DATA_TEMPR50[36] , 
        \R_DATA_TEMPR50[35] , \R_DATA_TEMPR50[34] , 
        \R_DATA_TEMPR50[33] , \R_DATA_TEMPR50[32] , 
        \R_DATA_TEMPR50[31] , \R_DATA_TEMPR50[30] , 
        \R_DATA_TEMPR50[29] , \R_DATA_TEMPR50[28] , 
        \R_DATA_TEMPR50[27] , \R_DATA_TEMPR50[26] , 
        \R_DATA_TEMPR50[25] , \R_DATA_TEMPR50[24] , 
        \R_DATA_TEMPR50[23] , \R_DATA_TEMPR50[22] , 
        \R_DATA_TEMPR50[21] , \R_DATA_TEMPR50[20] }), .B_DOUT({
        \R_DATA_TEMPR50[19] , \R_DATA_TEMPR50[18] , 
        \R_DATA_TEMPR50[17] , \R_DATA_TEMPR50[16] , 
        \R_DATA_TEMPR50[15] , \R_DATA_TEMPR50[14] , 
        \R_DATA_TEMPR50[13] , \R_DATA_TEMPR50[12] , 
        \R_DATA_TEMPR50[11] , \R_DATA_TEMPR50[10] , 
        \R_DATA_TEMPR50[9] , \R_DATA_TEMPR50[8] , \R_DATA_TEMPR50[7] , 
        \R_DATA_TEMPR50[6] , \R_DATA_TEMPR50[5] , \R_DATA_TEMPR50[4] , 
        \R_DATA_TEMPR50[3] , \R_DATA_TEMPR50[2] , \R_DATA_TEMPR50[1] , 
        \R_DATA_TEMPR50[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[50][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[12] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[12] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_239 (.A(\R_DATA_TEMPR24[30] ), .B(\R_DATA_TEMPR25[30] ), 
        .C(\R_DATA_TEMPR26[30] ), .D(\R_DATA_TEMPR27[30] ), .Y(
        OR4_239_Y));
    OR4 OR4_42 (.A(\R_DATA_TEMPR60[17] ), .B(\R_DATA_TEMPR61[17] ), .C(
        \R_DATA_TEMPR62[17] ), .D(\R_DATA_TEMPR63[17] ), .Y(OR4_42_Y));
    OR4 OR4_529 (.A(\R_DATA_TEMPR44[25] ), .B(\R_DATA_TEMPR45[25] ), 
        .C(\R_DATA_TEMPR46[25] ), .D(\R_DATA_TEMPR47[25] ), .Y(
        OR4_529_Y));
    OR4 OR4_477 (.A(\R_DATA_TEMPR28[28] ), .B(\R_DATA_TEMPR29[28] ), 
        .C(\R_DATA_TEMPR30[28] ), .D(\R_DATA_TEMPR31[28] ), .Y(
        OR4_477_Y));
    OR4 OR4_492 (.A(OR4_532_Y), .B(OR4_421_Y), .C(OR4_682_Y), .D(
        OR4_99_Y), .Y(OR4_492_Y));
    OR4 OR4_520 (.A(\R_DATA_TEMPR36[3] ), .B(\R_DATA_TEMPR37[3] ), .C(
        \R_DATA_TEMPR38[3] ), .D(\R_DATA_TEMPR39[3] ), .Y(OR4_520_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R59C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%59%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R59C0 (
        .A_DOUT({\R_DATA_TEMPR59[39] , \R_DATA_TEMPR59[38] , 
        \R_DATA_TEMPR59[37] , \R_DATA_TEMPR59[36] , 
        \R_DATA_TEMPR59[35] , \R_DATA_TEMPR59[34] , 
        \R_DATA_TEMPR59[33] , \R_DATA_TEMPR59[32] , 
        \R_DATA_TEMPR59[31] , \R_DATA_TEMPR59[30] , 
        \R_DATA_TEMPR59[29] , \R_DATA_TEMPR59[28] , 
        \R_DATA_TEMPR59[27] , \R_DATA_TEMPR59[26] , 
        \R_DATA_TEMPR59[25] , \R_DATA_TEMPR59[24] , 
        \R_DATA_TEMPR59[23] , \R_DATA_TEMPR59[22] , 
        \R_DATA_TEMPR59[21] , \R_DATA_TEMPR59[20] }), .B_DOUT({
        \R_DATA_TEMPR59[19] , \R_DATA_TEMPR59[18] , 
        \R_DATA_TEMPR59[17] , \R_DATA_TEMPR59[16] , 
        \R_DATA_TEMPR59[15] , \R_DATA_TEMPR59[14] , 
        \R_DATA_TEMPR59[13] , \R_DATA_TEMPR59[12] , 
        \R_DATA_TEMPR59[11] , \R_DATA_TEMPR59[10] , 
        \R_DATA_TEMPR59[9] , \R_DATA_TEMPR59[8] , \R_DATA_TEMPR59[7] , 
        \R_DATA_TEMPR59[6] , \R_DATA_TEMPR59[5] , \R_DATA_TEMPR59[4] , 
        \R_DATA_TEMPR59[3] , \R_DATA_TEMPR59[2] , \R_DATA_TEMPR59[1] , 
        \R_DATA_TEMPR59[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[59][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[14] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[14] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_499 (.A(\R_DATA_TEMPR12[27] ), .B(\R_DATA_TEMPR13[27] ), 
        .C(\R_DATA_TEMPR14[27] ), .D(\R_DATA_TEMPR15[27] ), .Y(
        OR4_499_Y));
    OR4 OR4_88 (.A(OR4_732_Y), .B(OR4_657_Y), .C(OR4_719_Y), .D(
        OR4_327_Y), .Y(OR4_88_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[7]  (.A(CFG3_15_Y), .B(CFG2_2_Y)
        , .Y(\BLKX2[7] ));
    OR4 OR4_205 (.A(\R_DATA_TEMPR44[26] ), .B(\R_DATA_TEMPR45[26] ), 
        .C(\R_DATA_TEMPR46[26] ), .D(\R_DATA_TEMPR47[26] ), .Y(
        OR4_205_Y));
    OR4 OR4_188 (.A(OR4_456_Y), .B(OR4_594_Y), .C(OR4_590_Y), .D(
        OR4_722_Y), .Y(OR4_188_Y));
    OR4 OR4_196 (.A(\R_DATA_TEMPR40[23] ), .B(\R_DATA_TEMPR41[23] ), 
        .C(\R_DATA_TEMPR42[23] ), .D(\R_DATA_TEMPR43[23] ), .Y(
        OR4_196_Y));
    OR4 OR4_112 (.A(\R_DATA_TEMPR32[33] ), .B(\R_DATA_TEMPR33[33] ), 
        .C(\R_DATA_TEMPR34[33] ), .D(\R_DATA_TEMPR35[33] ), .Y(
        OR4_112_Y));
    OR4 OR4_275 (.A(\R_DATA_TEMPR44[11] ), .B(\R_DATA_TEMPR45[11] ), 
        .C(\R_DATA_TEMPR46[11] ), .D(\R_DATA_TEMPR47[11] ), .Y(
        OR4_275_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R56C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%56%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R56C0 (
        .A_DOUT({\R_DATA_TEMPR56[39] , \R_DATA_TEMPR56[38] , 
        \R_DATA_TEMPR56[37] , \R_DATA_TEMPR56[36] , 
        \R_DATA_TEMPR56[35] , \R_DATA_TEMPR56[34] , 
        \R_DATA_TEMPR56[33] , \R_DATA_TEMPR56[32] , 
        \R_DATA_TEMPR56[31] , \R_DATA_TEMPR56[30] , 
        \R_DATA_TEMPR56[29] , \R_DATA_TEMPR56[28] , 
        \R_DATA_TEMPR56[27] , \R_DATA_TEMPR56[26] , 
        \R_DATA_TEMPR56[25] , \R_DATA_TEMPR56[24] , 
        \R_DATA_TEMPR56[23] , \R_DATA_TEMPR56[22] , 
        \R_DATA_TEMPR56[21] , \R_DATA_TEMPR56[20] }), .B_DOUT({
        \R_DATA_TEMPR56[19] , \R_DATA_TEMPR56[18] , 
        \R_DATA_TEMPR56[17] , \R_DATA_TEMPR56[16] , 
        \R_DATA_TEMPR56[15] , \R_DATA_TEMPR56[14] , 
        \R_DATA_TEMPR56[13] , \R_DATA_TEMPR56[12] , 
        \R_DATA_TEMPR56[11] , \R_DATA_TEMPR56[10] , 
        \R_DATA_TEMPR56[9] , \R_DATA_TEMPR56[8] , \R_DATA_TEMPR56[7] , 
        \R_DATA_TEMPR56[6] , \R_DATA_TEMPR56[5] , \R_DATA_TEMPR56[4] , 
        \R_DATA_TEMPR56[3] , \R_DATA_TEMPR56[2] , \R_DATA_TEMPR56[1] , 
        \R_DATA_TEMPR56[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[56][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[14] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[14] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_646 (.A(\R_DATA_TEMPR8[25] ), .B(\R_DATA_TEMPR9[25] ), .C(
        \R_DATA_TEMPR10[25] ), .D(\R_DATA_TEMPR11[25] ), .Y(OR4_646_Y));
    OR4 \OR4_R_DATA[37]  (.A(OR4_357_Y), .B(OR4_733_Y), .C(OR4_135_Y), 
        .D(OR4_218_Y), .Y(R_DATA[37]));
    OR4 OR4_257 (.A(\R_DATA_TEMPR20[14] ), .B(\R_DATA_TEMPR21[14] ), 
        .C(\R_DATA_TEMPR22[14] ), .D(\R_DATA_TEMPR23[14] ), .Y(
        OR4_257_Y));
    OR4 OR4_398 (.A(OR4_734_Y), .B(OR4_91_Y), .C(OR4_214_Y), .D(
        OR4_107_Y), .Y(OR4_398_Y));
    OR4 OR4_157 (.A(\R_DATA_TEMPR16[6] ), .B(\R_DATA_TEMPR17[6] ), .C(
        \R_DATA_TEMPR18[6] ), .D(\R_DATA_TEMPR19[6] ), .Y(OR4_157_Y));
    OR4 OR4_561 (.A(\R_DATA_TEMPR0[24] ), .B(\R_DATA_TEMPR1[24] ), .C(
        \R_DATA_TEMPR2[24] ), .D(\R_DATA_TEMPR3[24] ), .Y(OR4_561_Y));
    OR4 OR4_403 (.A(\R_DATA_TEMPR20[20] ), .B(\R_DATA_TEMPR21[20] ), 
        .C(\R_DATA_TEMPR22[20] ), .D(\R_DATA_TEMPR23[20] ), .Y(
        OR4_403_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R34C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%34%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R34C0 (
        .A_DOUT({\R_DATA_TEMPR34[39] , \R_DATA_TEMPR34[38] , 
        \R_DATA_TEMPR34[37] , \R_DATA_TEMPR34[36] , 
        \R_DATA_TEMPR34[35] , \R_DATA_TEMPR34[34] , 
        \R_DATA_TEMPR34[33] , \R_DATA_TEMPR34[32] , 
        \R_DATA_TEMPR34[31] , \R_DATA_TEMPR34[30] , 
        \R_DATA_TEMPR34[29] , \R_DATA_TEMPR34[28] , 
        \R_DATA_TEMPR34[27] , \R_DATA_TEMPR34[26] , 
        \R_DATA_TEMPR34[25] , \R_DATA_TEMPR34[24] , 
        \R_DATA_TEMPR34[23] , \R_DATA_TEMPR34[22] , 
        \R_DATA_TEMPR34[21] , \R_DATA_TEMPR34[20] }), .B_DOUT({
        \R_DATA_TEMPR34[19] , \R_DATA_TEMPR34[18] , 
        \R_DATA_TEMPR34[17] , \R_DATA_TEMPR34[16] , 
        \R_DATA_TEMPR34[15] , \R_DATA_TEMPR34[14] , 
        \R_DATA_TEMPR34[13] , \R_DATA_TEMPR34[12] , 
        \R_DATA_TEMPR34[11] , \R_DATA_TEMPR34[10] , 
        \R_DATA_TEMPR34[9] , \R_DATA_TEMPR34[8] , \R_DATA_TEMPR34[7] , 
        \R_DATA_TEMPR34[6] , \R_DATA_TEMPR34[5] , \R_DATA_TEMPR34[4] , 
        \R_DATA_TEMPR34[3] , \R_DATA_TEMPR34[2] , \R_DATA_TEMPR34[1] , 
        \R_DATA_TEMPR34[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[34][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[8] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[8] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_601 (.A(\R_DATA_TEMPR36[39] ), .B(\R_DATA_TEMPR37[39] ), 
        .C(\R_DATA_TEMPR38[39] ), .D(\R_DATA_TEMPR39[39] ), .Y(
        OR4_601_Y));
    CFG3 #( .INIT(8'h1) )  CFG3_7 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_7_Y));
    OR4 OR4_208 (.A(\R_DATA_TEMPR12[23] ), .B(\R_DATA_TEMPR13[23] ), 
        .C(\R_DATA_TEMPR14[23] ), .D(\R_DATA_TEMPR15[23] ), .Y(
        OR4_208_Y));
    OR4 OR4_219 (.A(\R_DATA_TEMPR16[12] ), .B(\R_DATA_TEMPR17[12] ), 
        .C(\R_DATA_TEMPR18[12] ), .D(\R_DATA_TEMPR19[12] ), .Y(
        OR4_219_Y));
    OR4 OR4_323 (.A(\R_DATA_TEMPR52[5] ), .B(\R_DATA_TEMPR53[5] ), .C(
        \R_DATA_TEMPR54[5] ), .D(\R_DATA_TEMPR55[5] ), .Y(OR4_323_Y));
    OR4 \OR4_R_DATA[19]  (.A(OR4_264_Y), .B(OR4_73_Y), .C(OR4_22_Y), 
        .D(OR4_686_Y), .Y(R_DATA[19]));
    OR4 OR4_720 (.A(\R_DATA_TEMPR36[36] ), .B(\R_DATA_TEMPR37[36] ), 
        .C(\R_DATA_TEMPR38[36] ), .D(\R_DATA_TEMPR39[36] ), .Y(
        OR4_720_Y));
    OR4 OR4_473 (.A(\R_DATA_TEMPR52[30] ), .B(\R_DATA_TEMPR53[30] ), 
        .C(\R_DATA_TEMPR54[30] ), .D(\R_DATA_TEMPR55[30] ), .Y(
        OR4_473_Y));
    OR4 OR4_671 (.A(\R_DATA_TEMPR40[4] ), .B(\R_DATA_TEMPR41[4] ), .C(
        \R_DATA_TEMPR42[4] ), .D(\R_DATA_TEMPR43[4] ), .Y(OR4_671_Y));
    OR4 OR4_737 (.A(\R_DATA_TEMPR8[32] ), .B(\R_DATA_TEMPR9[32] ), .C(
        \R_DATA_TEMPR10[32] ), .D(\R_DATA_TEMPR11[32] ), .Y(OR4_737_Y));
    OR4 OR4_422 (.A(\R_DATA_TEMPR0[37] ), .B(\R_DATA_TEMPR1[37] ), .C(
        \R_DATA_TEMPR2[37] ), .D(\R_DATA_TEMPR3[37] ), .Y(OR4_422_Y));
    OR4 OR4_278 (.A(\R_DATA_TEMPR44[38] ), .B(\R_DATA_TEMPR45[38] ), 
        .C(\R_DATA_TEMPR46[38] ), .D(\R_DATA_TEMPR47[38] ), .Y(
        OR4_278_Y));
    OR4 OR4_753 (.A(\R_DATA_TEMPR48[35] ), .B(\R_DATA_TEMPR49[35] ), 
        .C(\R_DATA_TEMPR50[35] ), .D(\R_DATA_TEMPR51[35] ), .Y(
        OR4_753_Y));
    OR4 OR4_734 (.A(\R_DATA_TEMPR32[10] ), .B(\R_DATA_TEMPR33[10] ), 
        .C(\R_DATA_TEMPR34[10] ), .D(\R_DATA_TEMPR35[10] ), .Y(
        OR4_734_Y));
    OR4 OR4_23 (.A(\R_DATA_TEMPR56[14] ), .B(\R_DATA_TEMPR57[14] ), .C(
        \R_DATA_TEMPR58[14] ), .D(\R_DATA_TEMPR59[14] ), .Y(OR4_23_Y));
    OR4 OR4_199 (.A(\R_DATA_TEMPR48[5] ), .B(\R_DATA_TEMPR49[5] ), .C(
        \R_DATA_TEMPR50[5] ), .D(\R_DATA_TEMPR51[5] ), .Y(OR4_199_Y));
    OR4 OR4_254 (.A(\R_DATA_TEMPR40[3] ), .B(\R_DATA_TEMPR41[3] ), .C(
        \R_DATA_TEMPR42[3] ), .D(\R_DATA_TEMPR43[3] ), .Y(OR4_254_Y));
    OR4 OR4_429 (.A(\R_DATA_TEMPR60[30] ), .B(\R_DATA_TEMPR61[30] ), 
        .C(\R_DATA_TEMPR62[30] ), .D(\R_DATA_TEMPR63[30] ), .Y(
        OR4_429_Y));
    OR4 OR4_262 (.A(\R_DATA_TEMPR40[15] ), .B(\R_DATA_TEMPR41[15] ), 
        .C(\R_DATA_TEMPR42[15] ), .D(\R_DATA_TEMPR43[15] ), .Y(
        OR4_262_Y));
    OR4 OR4_126 (.A(\R_DATA_TEMPR16[21] ), .B(\R_DATA_TEMPR17[21] ), 
        .C(\R_DATA_TEMPR18[21] ), .D(\R_DATA_TEMPR19[21] ), .Y(
        OR4_126_Y));
    OR4 OR4_94 (.A(\R_DATA_TEMPR12[20] ), .B(\R_DATA_TEMPR13[20] ), .C(
        \R_DATA_TEMPR14[20] ), .D(\R_DATA_TEMPR15[20] ), .Y(OR4_94_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%31%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R31C0 (
        .A_DOUT({\R_DATA_TEMPR31[39] , \R_DATA_TEMPR31[38] , 
        \R_DATA_TEMPR31[37] , \R_DATA_TEMPR31[36] , 
        \R_DATA_TEMPR31[35] , \R_DATA_TEMPR31[34] , 
        \R_DATA_TEMPR31[33] , \R_DATA_TEMPR31[32] , 
        \R_DATA_TEMPR31[31] , \R_DATA_TEMPR31[30] , 
        \R_DATA_TEMPR31[29] , \R_DATA_TEMPR31[28] , 
        \R_DATA_TEMPR31[27] , \R_DATA_TEMPR31[26] , 
        \R_DATA_TEMPR31[25] , \R_DATA_TEMPR31[24] , 
        \R_DATA_TEMPR31[23] , \R_DATA_TEMPR31[22] , 
        \R_DATA_TEMPR31[21] , \R_DATA_TEMPR31[20] }), .B_DOUT({
        \R_DATA_TEMPR31[19] , \R_DATA_TEMPR31[18] , 
        \R_DATA_TEMPR31[17] , \R_DATA_TEMPR31[16] , 
        \R_DATA_TEMPR31[15] , \R_DATA_TEMPR31[14] , 
        \R_DATA_TEMPR31[13] , \R_DATA_TEMPR31[12] , 
        \R_DATA_TEMPR31[11] , \R_DATA_TEMPR31[10] , 
        \R_DATA_TEMPR31[9] , \R_DATA_TEMPR31[8] , \R_DATA_TEMPR31[7] , 
        \R_DATA_TEMPR31[6] , \R_DATA_TEMPR31[5] , \R_DATA_TEMPR31[4] , 
        \R_DATA_TEMPR31[3] , \R_DATA_TEMPR31[2] , \R_DATA_TEMPR31[1] , 
        \R_DATA_TEMPR31[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[7] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[7] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_65 (.A(\R_DATA_TEMPR8[1] ), .B(\R_DATA_TEMPR9[1] ), .C(
        \R_DATA_TEMPR10[1] ), .D(\R_DATA_TEMPR11[1] ), .Y(OR4_65_Y));
    OR4 OR4_360 (.A(\R_DATA_TEMPR40[11] ), .B(\R_DATA_TEMPR41[11] ), 
        .C(\R_DATA_TEMPR42[11] ), .D(\R_DATA_TEMPR43[11] ), .Y(
        OR4_360_Y));
    OR4 OR4_355 (.A(\R_DATA_TEMPR60[31] ), .B(\R_DATA_TEMPR61[31] ), 
        .C(\R_DATA_TEMPR62[31] ), .D(\R_DATA_TEMPR63[31] ), .Y(
        OR4_355_Y));
    OR4 OR4_328 (.A(\R_DATA_TEMPR16[3] ), .B(\R_DATA_TEMPR17[3] ), .C(
        \R_DATA_TEMPR18[3] ), .D(\R_DATA_TEMPR19[3] ), .Y(OR4_328_Y));
    OR4 OR4_344 (.A(\R_DATA_TEMPR12[30] ), .B(\R_DATA_TEMPR13[30] ), 
        .C(\R_DATA_TEMPR14[30] ), .D(\R_DATA_TEMPR15[30] ), .Y(
        OR4_344_Y));
    OR4 OR4_185 (.A(\R_DATA_TEMPR8[17] ), .B(\R_DATA_TEMPR9[17] ), .C(
        \R_DATA_TEMPR10[17] ), .D(\R_DATA_TEMPR11[17] ), .Y(OR4_185_Y));
    OR4 OR4_141 (.A(OR4_14_Y), .B(OR4_181_Y), .C(OR4_280_Y), .D(
        OR4_51_Y), .Y(OR4_141_Y));
    OR4 OR4_717 (.A(\R_DATA_TEMPR24[2] ), .B(\R_DATA_TEMPR25[2] ), .C(
        \R_DATA_TEMPR26[2] ), .D(\R_DATA_TEMPR27[2] ), .Y(OR4_717_Y));
    OR4 OR4_36 (.A(OR4_783_Y), .B(OR4_606_Y), .C(OR4_791_Y), .D(
        OR4_344_Y), .Y(OR4_36_Y));
    OR4 OR4_487 (.A(\R_DATA_TEMPR32[20] ), .B(\R_DATA_TEMPR33[20] ), 
        .C(\R_DATA_TEMPR34[20] ), .D(\R_DATA_TEMPR35[20] ), .Y(
        OR4_487_Y));
    OR4 OR4_714 (.A(\R_DATA_TEMPR48[1] ), .B(\R_DATA_TEMPR49[1] ), .C(
        \R_DATA_TEMPR50[1] ), .D(\R_DATA_TEMPR51[1] ), .Y(OR4_714_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%22%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R22C0 (
        .A_DOUT({\R_DATA_TEMPR22[39] , \R_DATA_TEMPR22[38] , 
        \R_DATA_TEMPR22[37] , \R_DATA_TEMPR22[36] , 
        \R_DATA_TEMPR22[35] , \R_DATA_TEMPR22[34] , 
        \R_DATA_TEMPR22[33] , \R_DATA_TEMPR22[32] , 
        \R_DATA_TEMPR22[31] , \R_DATA_TEMPR22[30] , 
        \R_DATA_TEMPR22[29] , \R_DATA_TEMPR22[28] , 
        \R_DATA_TEMPR22[27] , \R_DATA_TEMPR22[26] , 
        \R_DATA_TEMPR22[25] , \R_DATA_TEMPR22[24] , 
        \R_DATA_TEMPR22[23] , \R_DATA_TEMPR22[22] , 
        \R_DATA_TEMPR22[21] , \R_DATA_TEMPR22[20] }), .B_DOUT({
        \R_DATA_TEMPR22[19] , \R_DATA_TEMPR22[18] , 
        \R_DATA_TEMPR22[17] , \R_DATA_TEMPR22[16] , 
        \R_DATA_TEMPR22[15] , \R_DATA_TEMPR22[14] , 
        \R_DATA_TEMPR22[13] , \R_DATA_TEMPR22[12] , 
        \R_DATA_TEMPR22[11] , \R_DATA_TEMPR22[10] , 
        \R_DATA_TEMPR22[9] , \R_DATA_TEMPR22[8] , \R_DATA_TEMPR22[7] , 
        \R_DATA_TEMPR22[6] , \R_DATA_TEMPR22[5] , \R_DATA_TEMPR22[4] , 
        \R_DATA_TEMPR22[3] , \R_DATA_TEMPR22[2] , \R_DATA_TEMPR22[1] , 
        \R_DATA_TEMPR22[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[5] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[5] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_501 (.A(OR4_34_Y), .B(OR4_186_Y), .C(OR4_716_Y), .D(
        OR4_335_Y), .Y(OR4_501_Y));
    OR4 OR4_21 (.A(\R_DATA_TEMPR48[34] ), .B(\R_DATA_TEMPR49[34] ), .C(
        \R_DATA_TEMPR50[34] ), .D(\R_DATA_TEMPR51[34] ), .Y(OR4_21_Y));
    OR4 OR4_129 (.A(\R_DATA_TEMPR16[13] ), .B(\R_DATA_TEMPR17[13] ), 
        .C(\R_DATA_TEMPR18[13] ), .D(\R_DATA_TEMPR19[13] ), .Y(
        OR4_129_Y));
    OR4 OR4_571 (.A(\R_DATA_TEMPR0[19] ), .B(\R_DATA_TEMPR1[19] ), .C(
        \R_DATA_TEMPR2[19] ), .D(\R_DATA_TEMPR3[19] ), .Y(OR4_571_Y));
    OR4 OR4_752 (.A(OR4_265_Y), .B(OR4_406_Y), .C(OR4_528_Y), .D(
        OR4_433_Y), .Y(OR4_752_Y));
    OR4 OR4_441 (.A(OR4_526_Y), .B(OR4_251_Y), .C(OR4_531_Y), .D(
        OR4_225_Y), .Y(OR4_441_Y));
    OR4 OR4_795 (.A(\R_DATA_TEMPR44[33] ), .B(\R_DATA_TEMPR45[33] ), 
        .C(\R_DATA_TEMPR46[33] ), .D(\R_DATA_TEMPR47[33] ), .Y(
        OR4_795_Y));
    OR4 OR4_697 (.A(OR4_215_Y), .B(OR4_677_Y), .C(OR4_709_Y), .D(
        OR4_316_Y), .Y(OR4_697_Y));
    OR4 OR4_448 (.A(\R_DATA_TEMPR24[17] ), .B(\R_DATA_TEMPR25[17] ), 
        .C(\R_DATA_TEMPR26[17] ), .D(\R_DATA_TEMPR27[17] ), .Y(
        OR4_448_Y));
    OR4 OR4_796 (.A(\R_DATA_TEMPR44[27] ), .B(\R_DATA_TEMPR45[27] ), 
        .C(\R_DATA_TEMPR46[27] ), .D(\R_DATA_TEMPR47[27] ), .Y(
        OR4_796_Y));
    OR4 OR4_285 (.A(OR4_718_Y), .B(OR4_473_Y), .C(OR4_496_Y), .D(
        OR4_429_Y), .Y(OR4_285_Y));
    OR4 OR4_202 (.A(\R_DATA_TEMPR36[18] ), .B(\R_DATA_TEMPR37[18] ), 
        .C(\R_DATA_TEMPR38[18] ), .D(\R_DATA_TEMPR39[18] ), .Y(
        OR4_202_Y));
    OR4 OR4_655 (.A(OR4_592_Y), .B(OR4_424_Y), .C(OR4_600_Y), .D(
        OR4_163_Y), .Y(OR4_655_Y));
    CFG3 #( .INIT(8'h80) )  CFG3_13 (.A(R_ADDR[13]), .B(R_ADDR[12]), 
        .C(R_ADDR[11]), .Y(CFG3_13_Y));
    OR4 OR4_272 (.A(\R_DATA_TEMPR52[21] ), .B(\R_DATA_TEMPR53[21] ), 
        .C(\R_DATA_TEMPR54[21] ), .D(\R_DATA_TEMPR55[21] ), .Y(
        OR4_272_Y));
    OR4 OR4_565 (.A(OR4_157_Y), .B(OR4_207_Y), .C(OR4_466_Y), .D(
        OR4_688_Y), .Y(OR4_565_Y));
    OR4 OR4_44 (.A(\R_DATA_TEMPR40[13] ), .B(\R_DATA_TEMPR41[13] ), .C(
        \R_DATA_TEMPR42[13] ), .D(\R_DATA_TEMPR43[13] ), .Y(OR4_44_Y));
    OR4 OR4_549 (.A(OR4_619_Y), .B(OR4_763_Y), .C(OR4_490_Y), .D(
        OR4_105_Y), .Y(OR4_549_Y));
    OR4 OR4_300 (.A(\R_DATA_TEMPR28[22] ), .B(\R_DATA_TEMPR29[22] ), 
        .C(\R_DATA_TEMPR30[22] ), .D(\R_DATA_TEMPR31[22] ), .Y(
        OR4_300_Y));
    OR4 OR4_435 (.A(\R_DATA_TEMPR36[9] ), .B(\R_DATA_TEMPR37[9] ), .C(
        \R_DATA_TEMPR38[9] ), .D(\R_DATA_TEMPR39[9] ), .Y(OR4_435_Y));
    OR4 OR4_540 (.A(\R_DATA_TEMPR16[2] ), .B(\R_DATA_TEMPR17[2] ), .C(
        \R_DATA_TEMPR18[2] ), .D(\R_DATA_TEMPR19[2] ), .Y(OR4_540_Y));
    OR4 OR4_483 (.A(OR4_374_Y), .B(OR4_715_Y), .C(OR4_178_Y), .D(
        OR4_683_Y), .Y(OR4_483_Y));
    OR4 OR4_681 (.A(\R_DATA_TEMPR44[36] ), .B(\R_DATA_TEMPR45[36] ), 
        .C(\R_DATA_TEMPR46[36] ), .D(\R_DATA_TEMPR47[36] ), .Y(
        OR4_681_Y));
    OR4 OR4_663 (.A(\R_DATA_TEMPR44[6] ), .B(\R_DATA_TEMPR45[6] ), .C(
        \R_DATA_TEMPR46[6] ), .D(\R_DATA_TEMPR47[6] ), .Y(OR4_663_Y));
    OR4 OR4_370 (.A(\R_DATA_TEMPR8[37] ), .B(\R_DATA_TEMPR9[37] ), .C(
        \R_DATA_TEMPR10[37] ), .D(\R_DATA_TEMPR11[37] ), .Y(OR4_370_Y));
    OR4 OR4_288 (.A(OR4_129_Y), .B(OR4_787_Y), .C(OR4_767_Y), .D(
        OR4_345_Y), .Y(OR4_288_Y));
    CFG3 #( .INIT(8'h4) )  CFG3_0 (.A(R_ADDR[13]), .B(R_ADDR[12]), .C(
        R_ADDR[11]), .Y(CFG3_0_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[8]  (.A(CFG3_10_Y), .B(CFG2_1_Y)
        , .Y(\BLKY2[8] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[12]  (.A(CFG3_3_Y), .B(CFG2_3_Y)
        , .Y(\BLKX2[12] ));
    OR4 OR4_30 (.A(OR4_362_Y), .B(OR4_511_Y), .C(OR4_249_Y), .D(
        OR4_663_Y), .Y(OR4_30_Y));
    OR4 OR4_650 (.A(\R_DATA_TEMPR12[29] ), .B(\R_DATA_TEMPR13[29] ), 
        .C(\R_DATA_TEMPR14[29] ), .D(\R_DATA_TEMPR15[29] ), .Y(
        OR4_650_Y));
    OR4 OR4_725 (.A(\R_DATA_TEMPR36[13] ), .B(\R_DATA_TEMPR37[13] ), 
        .C(\R_DATA_TEMPR38[13] ), .D(\R_DATA_TEMPR39[13] ), .Y(
        OR4_725_Y));
    OR4 OR4_627 (.A(OR4_213_Y), .B(OR4_118_Y), .C(OR4_631_Y), .D(
        OR4_79_Y), .Y(OR4_627_Y));
    OR4 OR4_297 (.A(\R_DATA_TEMPR56[27] ), .B(\R_DATA_TEMPR57[27] ), 
        .C(\R_DATA_TEMPR58[27] ), .D(\R_DATA_TEMPR59[27] ), .Y(
        OR4_297_Y));
    OR4 OR4_726 (.A(\R_DATA_TEMPR48[0] ), .B(\R_DATA_TEMPR49[0] ), .C(
        \R_DATA_TEMPR50[0] ), .D(\R_DATA_TEMPR51[0] ), .Y(OR4_726_Y));
    OR4 OR4_37 (.A(OR4_420_Y), .B(OR4_353_Y), .C(OR4_341_Y), .D(
        OR4_182_Y), .Y(OR4_37_Y));
    OR4 OR4_197 (.A(\R_DATA_TEMPR52[36] ), .B(\R_DATA_TEMPR53[36] ), 
        .C(\R_DATA_TEMPR54[36] ), .D(\R_DATA_TEMPR55[36] ), .Y(
        OR4_197_Y));
    OR4 OR4_357 (.A(OR4_422_Y), .B(OR4_53_Y), .C(OR4_370_Y), .D(
        OR4_745_Y), .Y(OR4_357_Y));
    OR4 OR4_150 (.A(\R_DATA_TEMPR16[35] ), .B(\R_DATA_TEMPR17[35] ), 
        .C(\R_DATA_TEMPR18[35] ), .D(\R_DATA_TEMPR19[35] ), .Y(
        OR4_150_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R43C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%43%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R43C0 (
        .A_DOUT({\R_DATA_TEMPR43[39] , \R_DATA_TEMPR43[38] , 
        \R_DATA_TEMPR43[37] , \R_DATA_TEMPR43[36] , 
        \R_DATA_TEMPR43[35] , \R_DATA_TEMPR43[34] , 
        \R_DATA_TEMPR43[33] , \R_DATA_TEMPR43[32] , 
        \R_DATA_TEMPR43[31] , \R_DATA_TEMPR43[30] , 
        \R_DATA_TEMPR43[29] , \R_DATA_TEMPR43[28] , 
        \R_DATA_TEMPR43[27] , \R_DATA_TEMPR43[26] , 
        \R_DATA_TEMPR43[25] , \R_DATA_TEMPR43[24] , 
        \R_DATA_TEMPR43[23] , \R_DATA_TEMPR43[22] , 
        \R_DATA_TEMPR43[21] , \R_DATA_TEMPR43[20] }), .B_DOUT({
        \R_DATA_TEMPR43[19] , \R_DATA_TEMPR43[18] , 
        \R_DATA_TEMPR43[17] , \R_DATA_TEMPR43[16] , 
        \R_DATA_TEMPR43[15] , \R_DATA_TEMPR43[14] , 
        \R_DATA_TEMPR43[13] , \R_DATA_TEMPR43[12] , 
        \R_DATA_TEMPR43[11] , \R_DATA_TEMPR43[10] , 
        \R_DATA_TEMPR43[9] , \R_DATA_TEMPR43[8] , \R_DATA_TEMPR43[7] , 
        \R_DATA_TEMPR43[6] , \R_DATA_TEMPR43[5] , \R_DATA_TEMPR43[4] , 
        \R_DATA_TEMPR43[3] , \R_DATA_TEMPR43[2] , \R_DATA_TEMPR43[1] , 
        \R_DATA_TEMPR43[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[43][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[10] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[10] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_434 (.A(\R_DATA_TEMPR60[3] ), .B(\R_DATA_TEMPR61[3] ), .C(
        \R_DATA_TEMPR62[3] ), .D(\R_DATA_TEMPR63[3] ), .Y(OR4_434_Y));
    OR4 OR4_163 (.A(\R_DATA_TEMPR12[10] ), .B(\R_DATA_TEMPR13[10] ), 
        .C(\R_DATA_TEMPR14[10] ), .D(\R_DATA_TEMPR15[10] ), .Y(
        OR4_163_Y));
    OR4 OR4_758 (.A(\R_DATA_TEMPR48[26] ), .B(\R_DATA_TEMPR49[26] ), 
        .C(\R_DATA_TEMPR50[26] ), .D(\R_DATA_TEMPR51[26] ), .Y(
        OR4_758_Y));
    OR4 OR4_343 (.A(\R_DATA_TEMPR12[32] ), .B(\R_DATA_TEMPR13[32] ), 
        .C(\R_DATA_TEMPR14[32] ), .D(\R_DATA_TEMPR15[32] ), .Y(
        OR4_343_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%10%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R10C0 (
        .A_DOUT({\R_DATA_TEMPR10[39] , \R_DATA_TEMPR10[38] , 
        \R_DATA_TEMPR10[37] , \R_DATA_TEMPR10[36] , 
        \R_DATA_TEMPR10[35] , \R_DATA_TEMPR10[34] , 
        \R_DATA_TEMPR10[33] , \R_DATA_TEMPR10[32] , 
        \R_DATA_TEMPR10[31] , \R_DATA_TEMPR10[30] , 
        \R_DATA_TEMPR10[29] , \R_DATA_TEMPR10[28] , 
        \R_DATA_TEMPR10[27] , \R_DATA_TEMPR10[26] , 
        \R_DATA_TEMPR10[25] , \R_DATA_TEMPR10[24] , 
        \R_DATA_TEMPR10[23] , \R_DATA_TEMPR10[22] , 
        \R_DATA_TEMPR10[21] , \R_DATA_TEMPR10[20] }), .B_DOUT({
        \R_DATA_TEMPR10[19] , \R_DATA_TEMPR10[18] , 
        \R_DATA_TEMPR10[17] , \R_DATA_TEMPR10[16] , 
        \R_DATA_TEMPR10[15] , \R_DATA_TEMPR10[14] , 
        \R_DATA_TEMPR10[13] , \R_DATA_TEMPR10[12] , 
        \R_DATA_TEMPR10[11] , \R_DATA_TEMPR10[10] , 
        \R_DATA_TEMPR10[9] , \R_DATA_TEMPR10[8] , \R_DATA_TEMPR10[7] , 
        \R_DATA_TEMPR10[6] , \R_DATA_TEMPR10[5] , \R_DATA_TEMPR10[4] , 
        \R_DATA_TEMPR10[3] , \R_DATA_TEMPR10[2] , \R_DATA_TEMPR10[1] , 
        \R_DATA_TEMPR10[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[2] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_740 (.A(\R_DATA_TEMPR60[7] ), .B(\R_DATA_TEMPR61[7] ), .C(
        \R_DATA_TEMPR62[7] ), .D(\R_DATA_TEMPR63[7] ), .Y(OR4_740_Y));
    OR4 OR4_336 (.A(\R_DATA_TEMPR48[19] ), .B(\R_DATA_TEMPR49[19] ), 
        .C(\R_DATA_TEMPR50[19] ), .D(\R_DATA_TEMPR51[19] ), .Y(
        OR4_336_Y));
    OR4 OR4_415 (.A(OR4_328_Y), .B(OR4_212_Y), .C(OR4_470_Y), .D(
        OR4_690_Y), .Y(OR4_415_Y));
    OR4 OR4_793 (.A(\R_DATA_TEMPR52[37] ), .B(\R_DATA_TEMPR53[37] ), 
        .C(\R_DATA_TEMPR54[37] ), .D(\R_DATA_TEMPR55[37] ), .Y(
        OR4_793_Y));
    OR4 OR4_442 (.A(OR4_756_Y), .B(OR4_232_Y), .C(OR4_567_Y), .D(
        OR4_96_Y), .Y(OR4_442_Y));
    OR4 OR4_294 (.A(\R_DATA_TEMPR32[30] ), .B(\R_DATA_TEMPR33[30] ), 
        .C(\R_DATA_TEMPR34[30] ), .D(\R_DATA_TEMPR35[30] ), .Y(
        OR4_294_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%19%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R19C0 (
        .A_DOUT({\R_DATA_TEMPR19[39] , \R_DATA_TEMPR19[38] , 
        \R_DATA_TEMPR19[37] , \R_DATA_TEMPR19[36] , 
        \R_DATA_TEMPR19[35] , \R_DATA_TEMPR19[34] , 
        \R_DATA_TEMPR19[33] , \R_DATA_TEMPR19[32] , 
        \R_DATA_TEMPR19[31] , \R_DATA_TEMPR19[30] , 
        \R_DATA_TEMPR19[29] , \R_DATA_TEMPR19[28] , 
        \R_DATA_TEMPR19[27] , \R_DATA_TEMPR19[26] , 
        \R_DATA_TEMPR19[25] , \R_DATA_TEMPR19[24] , 
        \R_DATA_TEMPR19[23] , \R_DATA_TEMPR19[22] , 
        \R_DATA_TEMPR19[21] , \R_DATA_TEMPR19[20] }), .B_DOUT({
        \R_DATA_TEMPR19[19] , \R_DATA_TEMPR19[18] , 
        \R_DATA_TEMPR19[17] , \R_DATA_TEMPR19[16] , 
        \R_DATA_TEMPR19[15] , \R_DATA_TEMPR19[14] , 
        \R_DATA_TEMPR19[13] , \R_DATA_TEMPR19[12] , 
        \R_DATA_TEMPR19[11] , \R_DATA_TEMPR19[10] , 
        \R_DATA_TEMPR19[9] , \R_DATA_TEMPR19[8] , \R_DATA_TEMPR19[7] , 
        \R_DATA_TEMPR19[6] , \R_DATA_TEMPR19[5] , \R_DATA_TEMPR19[4] , 
        \R_DATA_TEMPR19[3] , \R_DATA_TEMPR19[2] , \R_DATA_TEMPR19[1] , 
        \R_DATA_TEMPR19[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[4] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[4] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R52C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%52%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R52C0 (
        .A_DOUT({\R_DATA_TEMPR52[39] , \R_DATA_TEMPR52[38] , 
        \R_DATA_TEMPR52[37] , \R_DATA_TEMPR52[36] , 
        \R_DATA_TEMPR52[35] , \R_DATA_TEMPR52[34] , 
        \R_DATA_TEMPR52[33] , \R_DATA_TEMPR52[32] , 
        \R_DATA_TEMPR52[31] , \R_DATA_TEMPR52[30] , 
        \R_DATA_TEMPR52[29] , \R_DATA_TEMPR52[28] , 
        \R_DATA_TEMPR52[27] , \R_DATA_TEMPR52[26] , 
        \R_DATA_TEMPR52[25] , \R_DATA_TEMPR52[24] , 
        \R_DATA_TEMPR52[23] , \R_DATA_TEMPR52[22] , 
        \R_DATA_TEMPR52[21] , \R_DATA_TEMPR52[20] }), .B_DOUT({
        \R_DATA_TEMPR52[19] , \R_DATA_TEMPR52[18] , 
        \R_DATA_TEMPR52[17] , \R_DATA_TEMPR52[16] , 
        \R_DATA_TEMPR52[15] , \R_DATA_TEMPR52[14] , 
        \R_DATA_TEMPR52[13] , \R_DATA_TEMPR52[12] , 
        \R_DATA_TEMPR52[11] , \R_DATA_TEMPR52[10] , 
        \R_DATA_TEMPR52[9] , \R_DATA_TEMPR52[8] , \R_DATA_TEMPR52[7] , 
        \R_DATA_TEMPR52[6] , \R_DATA_TEMPR52[5] , \R_DATA_TEMPR52[4] , 
        \R_DATA_TEMPR52[3] , \R_DATA_TEMPR52[2] , \R_DATA_TEMPR52[1] , 
        \R_DATA_TEMPR52[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[52][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[13] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[13] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_449 (.A(\R_DATA_TEMPR0[28] ), .B(\R_DATA_TEMPR1[28] ), .C(
        \R_DATA_TEMPR2[28] ), .D(\R_DATA_TEMPR3[28] ), .Y(OR4_449_Y));
    OR4 OR4_505 (.A(\R_DATA_TEMPR20[28] ), .B(\R_DATA_TEMPR21[28] ), 
        .C(\R_DATA_TEMPR22[28] ), .D(\R_DATA_TEMPR23[28] ), .Y(
        OR4_505_Y));
    OR4 \OR4_R_DATA[24]  (.A(OR4_692_Y), .B(OR4_417_Y), .C(OR4_5_Y), 
        .D(OR4_356_Y), .Y(R_DATA[24]));
    OR4 OR4_85 (.A(\R_DATA_TEMPR32[29] ), .B(\R_DATA_TEMPR33[29] ), .C(
        \R_DATA_TEMPR34[29] ), .D(\R_DATA_TEMPR35[29] ), .Y(OR4_85_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%5%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R5C0 (.A_DOUT({
        \R_DATA_TEMPR5[39] , \R_DATA_TEMPR5[38] , \R_DATA_TEMPR5[37] , 
        \R_DATA_TEMPR5[36] , \R_DATA_TEMPR5[35] , \R_DATA_TEMPR5[34] , 
        \R_DATA_TEMPR5[33] , \R_DATA_TEMPR5[32] , \R_DATA_TEMPR5[31] , 
        \R_DATA_TEMPR5[30] , \R_DATA_TEMPR5[29] , \R_DATA_TEMPR5[28] , 
        \R_DATA_TEMPR5[27] , \R_DATA_TEMPR5[26] , \R_DATA_TEMPR5[25] , 
        \R_DATA_TEMPR5[24] , \R_DATA_TEMPR5[23] , \R_DATA_TEMPR5[22] , 
        \R_DATA_TEMPR5[21] , \R_DATA_TEMPR5[20] }), .B_DOUT({
        \R_DATA_TEMPR5[19] , \R_DATA_TEMPR5[18] , \R_DATA_TEMPR5[17] , 
        \R_DATA_TEMPR5[16] , \R_DATA_TEMPR5[15] , \R_DATA_TEMPR5[14] , 
        \R_DATA_TEMPR5[13] , \R_DATA_TEMPR5[12] , \R_DATA_TEMPR5[11] , 
        \R_DATA_TEMPR5[10] , \R_DATA_TEMPR5[9] , \R_DATA_TEMPR5[8] , 
        \R_DATA_TEMPR5[7] , \R_DATA_TEMPR5[6] , \R_DATA_TEMPR5[5] , 
        \R_DATA_TEMPR5[4] , \R_DATA_TEMPR5[3] , \R_DATA_TEMPR5[2] , 
        \R_DATA_TEMPR5[1] , \R_DATA_TEMPR5[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[5][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_146 (.A(OR4_380_Y), .B(OR4_390_Y), .C(OR4_381_Y), .D(
        OR4_233_Y), .Y(OR4_146_Y));
    OR4 OR4_158 (.A(\R_DATA_TEMPR24[32] ), .B(\R_DATA_TEMPR25[32] ), 
        .C(\R_DATA_TEMPR26[32] ), .D(\R_DATA_TEMPR27[32] ), .Y(
        OR4_158_Y));
    OR4 \OR4_R_DATA[12]  (.A(OR4_573_Y), .B(OR4_554_Y), .C(OR4_446_Y), 
        .D(OR4_80_Y), .Y(R_DATA[12]));
    CFG3 #( .INIT(8'h1) )  CFG3_10 (.A(R_ADDR[13]), .B(R_ADDR[12]), .C(
        R_ADDR[11]), .Y(CFG3_10_Y));
    OR4 OR4_581 (.A(OR4_294_Y), .B(OR4_203_Y), .C(OR4_707_Y), .D(
        OR4_161_Y), .Y(OR4_581_Y));
    OR4 OR4_575 (.A(\R_DATA_TEMPR52[12] ), .B(\R_DATA_TEMPR53[12] ), 
        .C(\R_DATA_TEMPR54[12] ), .D(\R_DATA_TEMPR55[12] ), .Y(
        OR4_575_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%16%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R16C0 (
        .A_DOUT({\R_DATA_TEMPR16[39] , \R_DATA_TEMPR16[38] , 
        \R_DATA_TEMPR16[37] , \R_DATA_TEMPR16[36] , 
        \R_DATA_TEMPR16[35] , \R_DATA_TEMPR16[34] , 
        \R_DATA_TEMPR16[33] , \R_DATA_TEMPR16[32] , 
        \R_DATA_TEMPR16[31] , \R_DATA_TEMPR16[30] , 
        \R_DATA_TEMPR16[29] , \R_DATA_TEMPR16[28] , 
        \R_DATA_TEMPR16[27] , \R_DATA_TEMPR16[26] , 
        \R_DATA_TEMPR16[25] , \R_DATA_TEMPR16[24] , 
        \R_DATA_TEMPR16[23] , \R_DATA_TEMPR16[22] , 
        \R_DATA_TEMPR16[21] , \R_DATA_TEMPR16[20] }), .B_DOUT({
        \R_DATA_TEMPR16[19] , \R_DATA_TEMPR16[18] , 
        \R_DATA_TEMPR16[17] , \R_DATA_TEMPR16[16] , 
        \R_DATA_TEMPR16[15] , \R_DATA_TEMPR16[14] , 
        \R_DATA_TEMPR16[13] , \R_DATA_TEMPR16[12] , 
        \R_DATA_TEMPR16[11] , \R_DATA_TEMPR16[10] , 
        \R_DATA_TEMPR16[9] , \R_DATA_TEMPR16[8] , \R_DATA_TEMPR16[7] , 
        \R_DATA_TEMPR16[6] , \R_DATA_TEMPR16[5] , \R_DATA_TEMPR16[4] , 
        \R_DATA_TEMPR16[3] , \R_DATA_TEMPR16[2] , \R_DATA_TEMPR16[1] , 
        \R_DATA_TEMPR16[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[4] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_603 (.A(OR4_21_Y), .B(OR4_574_Y), .C(OR4_605_Y), .D(
        OR4_61_Y), .Y(OR4_603_Y));
    OR4 OR4_69 (.A(\R_DATA_TEMPR20[33] ), .B(\R_DATA_TEMPR21[33] ), .C(
        \R_DATA_TEMPR22[33] ), .D(\R_DATA_TEMPR23[33] ), .Y(OR4_69_Y));
    OR4 OR4_227 (.A(\R_DATA_TEMPR52[28] ), .B(\R_DATA_TEMPR53[28] ), 
        .C(\R_DATA_TEMPR54[28] ), .D(\R_DATA_TEMPR55[28] ), .Y(
        OR4_227_Y));
    OR4 OR4_673 (.A(\R_DATA_TEMPR60[33] ), .B(\R_DATA_TEMPR61[33] ), 
        .C(\R_DATA_TEMPR62[33] ), .D(\R_DATA_TEMPR63[33] ), .Y(
        OR4_673_Y));
    OR4 OR4_395 (.A(\R_DATA_TEMPR60[36] ), .B(\R_DATA_TEMPR61[36] ), 
        .C(\R_DATA_TEMPR62[36] ), .D(\R_DATA_TEMPR63[36] ), .Y(
        OR4_395_Y));
    OR4 OR4_414 (.A(\R_DATA_TEMPR56[5] ), .B(\R_DATA_TEMPR57[5] ), .C(
        \R_DATA_TEMPR58[5] ), .D(\R_DATA_TEMPR59[5] ), .Y(OR4_414_Y));
    OR4 OR4_127 (.A(\R_DATA_TEMPR36[15] ), .B(\R_DATA_TEMPR37[15] ), 
        .C(\R_DATA_TEMPR38[15] ), .D(\R_DATA_TEMPR39[15] ), .Y(
        OR4_127_Y));
    OR4 OR4_348 (.A(\R_DATA_TEMPR36[31] ), .B(\R_DATA_TEMPR37[31] ), 
        .C(\R_DATA_TEMPR38[31] ), .D(\R_DATA_TEMPR39[31] ), .Y(
        OR4_348_Y));
    OR4 OR4_162 (.A(\R_DATA_TEMPR12[12] ), .B(\R_DATA_TEMPR13[12] ), 
        .C(\R_DATA_TEMPR14[12] ), .D(\R_DATA_TEMPR15[12] ), .Y(
        OR4_162_Y));
    OR4 OR4_282 (.A(\R_DATA_TEMPR60[9] ), .B(\R_DATA_TEMPR61[9] ), .C(
        \R_DATA_TEMPR62[9] ), .D(\R_DATA_TEMPR63[9] ), .Y(OR4_282_Y));
    OR4 OR4_316 (.A(\R_DATA_TEMPR12[15] ), .B(\R_DATA_TEMPR13[15] ), 
        .C(\R_DATA_TEMPR14[15] ), .D(\R_DATA_TEMPR15[15] ), .Y(
        OR4_316_Y));
    OR4 OR4_134 (.A(OR4_261_Y), .B(OR4_379_Y), .C(OR4_469_Y), .D(
        OR4_584_Y), .Y(OR4_134_Y));
    OR4 OR4_723 (.A(\R_DATA_TEMPR0[12] ), .B(\R_DATA_TEMPR1[12] ), .C(
        \R_DATA_TEMPR2[12] ), .D(\R_DATA_TEMPR3[12] ), .Y(OR4_723_Y));
    OR4 OR4_103 (.A(\R_DATA_TEMPR0[6] ), .B(\R_DATA_TEMPR1[6] ), .C(
        \R_DATA_TEMPR2[6] ), .D(\R_DATA_TEMPR3[6] ), .Y(OR4_103_Y));
    OR4 OR4_224 (.A(OR4_338_Y), .B(OR4_252_Y), .C(OR4_239_Y), .D(
        OR4_70_Y), .Y(OR4_224_Y));
    OR4 OR4_149 (.A(OR4_457_Y), .B(OR4_616_Y), .C(OR4_727_Y), .D(
        OR4_641_Y), .Y(OR4_149_Y));
    OR4 OR4_792 (.A(\R_DATA_TEMPR32[4] ), .B(\R_DATA_TEMPR33[4] ), .C(
        \R_DATA_TEMPR34[4] ), .D(\R_DATA_TEMPR35[4] ), .Y(OR4_792_Y));
    OR4 OR4_380 (.A(\R_DATA_TEMPR16[31] ), .B(\R_DATA_TEMPR17[31] ), 
        .C(\R_DATA_TEMPR18[31] ), .D(\R_DATA_TEMPR19[31] ), .Y(
        OR4_380_Y));
    OR4 \OR4_R_DATA[13]  (.A(OR4_484_Y), .B(OR4_288_Y), .C(OR4_255_Y), 
        .D(OR4_231_Y), .Y(R_DATA[13]));
    OR4 OR4_173 (.A(\R_DATA_TEMPR24[15] ), .B(\R_DATA_TEMPR25[15] ), 
        .C(\R_DATA_TEMPR26[15] ), .D(\R_DATA_TEMPR27[15] ), .Y(
        OR4_173_Y));
    OR4 OR4_269 (.A(\R_DATA_TEMPR12[18] ), .B(\R_DATA_TEMPR13[18] ), 
        .C(\R_DATA_TEMPR14[18] ), .D(\R_DATA_TEMPR15[18] ), .Y(
        OR4_269_Y));
    OR4 OR4_731 (.A(OR4_209_Y), .B(OR4_342_Y), .C(OR4_340_Y), .D(
        OR4_471_Y), .Y(OR4_731_Y));
    OR4 OR4_695 (.A(\R_DATA_TEMPR36[22] ), .B(\R_DATA_TEMPR37[22] ), 
        .C(\R_DATA_TEMPR38[22] ), .D(\R_DATA_TEMPR39[22] ), .Y(
        OR4_695_Y));
    OR4 OR4_62 (.A(OR4_45_Y), .B(OR4_200_Y), .C(OR4_317_Y), .D(
        OR4_228_Y), .Y(OR4_62_Y));
    OR4 OR4_38 (.A(\R_DATA_TEMPR52[1] ), .B(\R_DATA_TEMPR53[1] ), .C(
        \R_DATA_TEMPR54[1] ), .D(\R_DATA_TEMPR55[1] ), .Y(OR4_38_Y));
    OR4 OR4_325 (.A(\R_DATA_TEMPR32[23] ), .B(\R_DATA_TEMPR33[23] ), 
        .C(\R_DATA_TEMPR34[23] ), .D(\R_DATA_TEMPR35[23] ), .Y(
        OR4_325_Y));
    OR4 OR4_536 (.A(\R_DATA_TEMPR32[25] ), .B(\R_DATA_TEMPR33[25] ), 
        .C(\R_DATA_TEMPR34[25] ), .D(\R_DATA_TEMPR35[25] ), .Y(
        OR4_536_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R48C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%48%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R48C0 (
        .A_DOUT({\R_DATA_TEMPR48[39] , \R_DATA_TEMPR48[38] , 
        \R_DATA_TEMPR48[37] , \R_DATA_TEMPR48[36] , 
        \R_DATA_TEMPR48[35] , \R_DATA_TEMPR48[34] , 
        \R_DATA_TEMPR48[33] , \R_DATA_TEMPR48[32] , 
        \R_DATA_TEMPR48[31] , \R_DATA_TEMPR48[30] , 
        \R_DATA_TEMPR48[29] , \R_DATA_TEMPR48[28] , 
        \R_DATA_TEMPR48[27] , \R_DATA_TEMPR48[26] , 
        \R_DATA_TEMPR48[25] , \R_DATA_TEMPR48[24] , 
        \R_DATA_TEMPR48[23] , \R_DATA_TEMPR48[22] , 
        \R_DATA_TEMPR48[21] , \R_DATA_TEMPR48[20] }), .B_DOUT({
        \R_DATA_TEMPR48[19] , \R_DATA_TEMPR48[18] , 
        \R_DATA_TEMPR48[17] , \R_DATA_TEMPR48[16] , 
        \R_DATA_TEMPR48[15] , \R_DATA_TEMPR48[14] , 
        \R_DATA_TEMPR48[13] , \R_DATA_TEMPR48[12] , 
        \R_DATA_TEMPR48[11] , \R_DATA_TEMPR48[10] , 
        \R_DATA_TEMPR48[9] , \R_DATA_TEMPR48[8] , \R_DATA_TEMPR48[7] , 
        \R_DATA_TEMPR48[6] , \R_DATA_TEMPR48[5] , \R_DATA_TEMPR48[4] , 
        \R_DATA_TEMPR48[3] , \R_DATA_TEMPR48[2] , \R_DATA_TEMPR48[1] , 
        \R_DATA_TEMPR48[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[48][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[12] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[12] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_114 (.A(\R_DATA_TEMPR0[8] ), .B(\R_DATA_TEMPR1[8] ), .C(
        \R_DATA_TEMPR2[8] ), .D(\R_DATA_TEMPR3[8] ), .Y(OR4_114_Y));
    OR4 OR4_155 (.A(OR4_66_Y), .B(OR4_742_Y), .C(OR4_612_Y), .D(
        OR4_26_Y), .Y(OR4_155_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[6]  (.A(CFG3_5_Y), .B(CFG2_2_Y), 
        .Y(\BLKX2[6] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[14]  (.A(CFG3_5_Y), .B(CFG2_3_Y)
        , .Y(\BLKX2[14] ));
    OR4 OR4_457 (.A(\R_DATA_TEMPR32[16] ), .B(\R_DATA_TEMPR33[16] ), 
        .C(\R_DATA_TEMPR34[16] ), .D(\R_DATA_TEMPR35[16] ), .Y(
        OR4_457_Y));
    OR4 OR4_102 (.A(\R_DATA_TEMPR0[32] ), .B(\R_DATA_TEMPR1[32] ), .C(
        \R_DATA_TEMPR2[32] ), .D(\R_DATA_TEMPR3[32] ), .Y(OR4_102_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%25%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R25C0 (
        .A_DOUT({\R_DATA_TEMPR25[39] , \R_DATA_TEMPR25[38] , 
        \R_DATA_TEMPR25[37] , \R_DATA_TEMPR25[36] , 
        \R_DATA_TEMPR25[35] , \R_DATA_TEMPR25[34] , 
        \R_DATA_TEMPR25[33] , \R_DATA_TEMPR25[32] , 
        \R_DATA_TEMPR25[31] , \R_DATA_TEMPR25[30] , 
        \R_DATA_TEMPR25[29] , \R_DATA_TEMPR25[28] , 
        \R_DATA_TEMPR25[27] , \R_DATA_TEMPR25[26] , 
        \R_DATA_TEMPR25[25] , \R_DATA_TEMPR25[24] , 
        \R_DATA_TEMPR25[23] , \R_DATA_TEMPR25[22] , 
        \R_DATA_TEMPR25[21] , \R_DATA_TEMPR25[20] }), .B_DOUT({
        \R_DATA_TEMPR25[19] , \R_DATA_TEMPR25[18] , 
        \R_DATA_TEMPR25[17] , \R_DATA_TEMPR25[16] , 
        \R_DATA_TEMPR25[15] , \R_DATA_TEMPR25[14] , 
        \R_DATA_TEMPR25[13] , \R_DATA_TEMPR25[12] , 
        \R_DATA_TEMPR25[11] , \R_DATA_TEMPR25[10] , 
        \R_DATA_TEMPR25[9] , \R_DATA_TEMPR25[8] , \R_DATA_TEMPR25[7] , 
        \R_DATA_TEMPR25[6] , \R_DATA_TEMPR25[5] , \R_DATA_TEMPR25[4] , 
        \R_DATA_TEMPR25[3] , \R_DATA_TEMPR25[2] , \R_DATA_TEMPR25[1] , 
        \R_DATA_TEMPR25[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[6] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    CFG1 #( .INIT(2'h1) )  \INVBLKY0[0]  (.A(R_ADDR[9]), .Y(\BLKY0[0] )
        );
    OR4 OR4_690 (.A(\R_DATA_TEMPR28[3] ), .B(\R_DATA_TEMPR29[3] ), .C(
        \R_DATA_TEMPR30[3] ), .D(\R_DATA_TEMPR31[3] ), .Y(OR4_690_Y));
    OR4 OR4_722 (.A(\R_DATA_TEMPR12[31] ), .B(\R_DATA_TEMPR13[31] ), 
        .C(\R_DATA_TEMPR14[31] ), .D(\R_DATA_TEMPR15[31] ), .Y(
        OR4_722_Y));
    OR4 OR4_172 (.A(\R_DATA_TEMPR52[17] ), .B(\R_DATA_TEMPR53[17] ), 
        .C(\R_DATA_TEMPR54[17] ), .D(\R_DATA_TEMPR55[17] ), .Y(
        OR4_172_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R60C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%60%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R60C0 (
        .A_DOUT({\R_DATA_TEMPR60[39] , \R_DATA_TEMPR60[38] , 
        \R_DATA_TEMPR60[37] , \R_DATA_TEMPR60[36] , 
        \R_DATA_TEMPR60[35] , \R_DATA_TEMPR60[34] , 
        \R_DATA_TEMPR60[33] , \R_DATA_TEMPR60[32] , 
        \R_DATA_TEMPR60[31] , \R_DATA_TEMPR60[30] , 
        \R_DATA_TEMPR60[29] , \R_DATA_TEMPR60[28] , 
        \R_DATA_TEMPR60[27] , \R_DATA_TEMPR60[26] , 
        \R_DATA_TEMPR60[25] , \R_DATA_TEMPR60[24] , 
        \R_DATA_TEMPR60[23] , \R_DATA_TEMPR60[22] , 
        \R_DATA_TEMPR60[21] , \R_DATA_TEMPR60[20] }), .B_DOUT({
        \R_DATA_TEMPR60[19] , \R_DATA_TEMPR60[18] , 
        \R_DATA_TEMPR60[17] , \R_DATA_TEMPR60[16] , 
        \R_DATA_TEMPR60[15] , \R_DATA_TEMPR60[14] , 
        \R_DATA_TEMPR60[13] , \R_DATA_TEMPR60[12] , 
        \R_DATA_TEMPR60[11] , \R_DATA_TEMPR60[10] , 
        \R_DATA_TEMPR60[9] , \R_DATA_TEMPR60[8] , \R_DATA_TEMPR60[7] , 
        \R_DATA_TEMPR60[6] , \R_DATA_TEMPR60[5] , \R_DATA_TEMPR60[4] , 
        \R_DATA_TEMPR60[3] , \R_DATA_TEMPR60[2] , \R_DATA_TEMPR60[1] , 
        \R_DATA_TEMPR60[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[60][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[15] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[15] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_745 (.A(\R_DATA_TEMPR12[37] ), .B(\R_DATA_TEMPR13[37] ), 
        .C(\R_DATA_TEMPR14[37] ), .D(\R_DATA_TEMPR15[37] ), .Y(
        OR4_745_Y));
    OR4 OR4_647 (.A(\R_DATA_TEMPR56[12] ), .B(\R_DATA_TEMPR57[12] ), 
        .C(\R_DATA_TEMPR58[12] ), .D(\R_DATA_TEMPR59[12] ), .Y(
        OR4_647_Y));
    OR4 OR4_746 (.A(\R_DATA_TEMPR56[7] ), .B(\R_DATA_TEMPR57[7] ), .C(
        \R_DATA_TEMPR58[7] ), .D(\R_DATA_TEMPR59[7] ), .Y(OR4_746_Y));
    OR4 OR4_711 (.A(\R_DATA_TEMPR28[33] ), .B(\R_DATA_TEMPR29[33] ), 
        .C(\R_DATA_TEMPR30[33] ), .D(\R_DATA_TEMPR31[33] ), .Y(
        OR4_711_Y));
    OR4 OR4_585 (.A(OR4_527_Y), .B(OR4_358_Y), .C(OR4_537_Y), .D(
        OR4_94_Y), .Y(OR4_585_Y));
    OR4 OR4_767 (.A(\R_DATA_TEMPR24[13] ), .B(\R_DATA_TEMPR25[13] ), 
        .C(\R_DATA_TEMPR26[13] ), .D(\R_DATA_TEMPR27[13] ), .Y(
        OR4_767_Y));
    OR4 OR4_255 (.A(OR4_569_Y), .B(OR4_725_Y), .C(OR4_44_Y), .D(
        OR4_744_Y), .Y(OR4_255_Y));
    OR4 OR4_397 (.A(OR4_540_Y), .B(OR4_450_Y), .C(OR4_717_Y), .D(
        OR4_132_Y), .Y(OR4_397_Y));
    OR4 OR4_190 (.A(\R_DATA_TEMPR12[28] ), .B(\R_DATA_TEMPR13[28] ), 
        .C(\R_DATA_TEMPR14[28] ), .D(\R_DATA_TEMPR15[28] ), .Y(
        OR4_190_Y));
    OR4 OR4_764 (.A(\R_DATA_TEMPR52[18] ), .B(\R_DATA_TEMPR53[18] ), 
        .C(\R_DATA_TEMPR54[18] ), .D(\R_DATA_TEMPR55[18] ), .Y(
        OR4_764_Y));
    OR4 OR4_625 (.A(\R_DATA_TEMPR16[37] ), .B(\R_DATA_TEMPR17[37] ), 
        .C(\R_DATA_TEMPR18[37] ), .D(\R_DATA_TEMPR19[37] ), .Y(
        OR4_625_Y));
    OR4 OR4_538 (.A(\R_DATA_TEMPR48[7] ), .B(\R_DATA_TEMPR49[7] ), .C(
        \R_DATA_TEMPR50[7] ), .D(\R_DATA_TEMPR51[7] ), .Y(OR4_538_Y));
    OR4 OR4_26 (.A(\R_DATA_TEMPR60[23] ), .B(\R_DATA_TEMPR61[23] ), .C(
        \R_DATA_TEMPR62[23] ), .D(\R_DATA_TEMPR63[23] ), .Y(OR4_26_Y));
    OR4 OR4_53 (.A(\R_DATA_TEMPR4[37] ), .B(\R_DATA_TEMPR5[37] ), .C(
        \R_DATA_TEMPR6[37] ), .D(\R_DATA_TEMPR7[37] ), .Y(OR4_53_Y));
    OR4 OR4_683 (.A(\R_DATA_TEMPR28[27] ), .B(\R_DATA_TEMPR29[27] ), 
        .C(\R_DATA_TEMPR30[27] ), .D(\R_DATA_TEMPR31[27] ), .Y(
        OR4_683_Y));
    OR4 OR4_209 (.A(\R_DATA_TEMPR0[21] ), .B(\R_DATA_TEMPR1[21] ), .C(
        \R_DATA_TEMPR2[21] ), .D(\R_DATA_TEMPR3[21] ), .Y(OR4_209_Y));
    OR4 OR4_798 (.A(\R_DATA_TEMPR4[14] ), .B(\R_DATA_TEMPR5[14] ), .C(
        \R_DATA_TEMPR6[14] ), .D(\R_DATA_TEMPR7[14] ), .Y(OR4_798_Y));
    OR4 OR4_516 (.A(\R_DATA_TEMPR36[37] ), .B(\R_DATA_TEMPR37[37] ), 
        .C(\R_DATA_TEMPR38[37] ), .D(\R_DATA_TEMPR39[37] ), .Y(
        OR4_516_Y));
    OR4 OR4_279 (.A(OR4_644_Y), .B(OR4_396_Y), .C(OR4_427_Y), .D(
        OR4_145_Y), .Y(OR4_279_Y));
    OR4 OR4_436 (.A(OR4_112_Y), .B(OR4_32_Y), .C(OR4_542_Y), .D(
        OR4_795_Y), .Y(OR4_436_Y));
    OR4 OR4_89 (.A(\R_DATA_TEMPR24[4] ), .B(\R_DATA_TEMPR25[4] ), .C(
        \R_DATA_TEMPR26[4] ), .D(\R_DATA_TEMPR27[4] ), .Y(OR4_89_Y));
    OR4 OR4_453 (.A(\R_DATA_TEMPR12[33] ), .B(\R_DATA_TEMPR13[33] ), 
        .C(\R_DATA_TEMPR14[33] ), .D(\R_DATA_TEMPR15[33] ), .Y(
        OR4_453_Y));
    OR4 OR4_651 (.A(\R_DATA_TEMPR56[31] ), .B(\R_DATA_TEMPR57[31] ), 
        .C(\R_DATA_TEMPR58[31] ), .D(\R_DATA_TEMPR59[31] ), .Y(
        OR4_651_Y));
    OR4 OR4_198 (.A(\R_DATA_TEMPR16[16] ), .B(\R_DATA_TEMPR17[16] ), 
        .C(\R_DATA_TEMPR18[16] ), .D(\R_DATA_TEMPR19[16] ), .Y(
        OR4_198_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[3]  (.A(CFG3_2_Y), .B(CFG2_2_Y), 
        .Y(\BLKX2[3] ));
    OR4 OR4_258 (.A(\R_DATA_TEMPR20[18] ), .B(\R_DATA_TEMPR21[18] ), 
        .C(\R_DATA_TEMPR22[18] ), .D(\R_DATA_TEMPR23[18] ), .Y(
        OR4_258_Y));
    OR4 \OR4_R_DATA[21]  (.A(OR4_731_Y), .B(OR4_696_Y), .C(OR4_710_Y), 
        .D(OR4_459_Y), .Y(R_DATA[21]));
    OR4 OR4_620 (.A(OR4_175_Y), .B(OR4_304_Y), .C(OR4_386_Y), .D(
        OR4_282_Y), .Y(OR4_620_Y));
    OR4 OR4_183 (.A(\R_DATA_TEMPR40[5] ), .B(\R_DATA_TEMPR41[5] ), .C(
        \R_DATA_TEMPR42[5] ), .D(\R_DATA_TEMPR43[5] ), .Y(OR4_183_Y));
    OR4 OR4_332 (.A(OR4_4_Y), .B(OR4_720_Y), .C(OR4_428_Y), .D(
        OR4_681_Y), .Y(OR4_332_Y));
    OR4 OR4_13 (.A(\R_DATA_TEMPR24[21] ), .B(\R_DATA_TEMPR25[21] ), .C(
        \R_DATA_TEMPR26[21] ), .D(\R_DATA_TEMPR27[21] ), .Y(OR4_13_Y));
    OR4 OR4_247 (.A(\R_DATA_TEMPR12[5] ), .B(\R_DATA_TEMPR13[5] ), .C(
        \R_DATA_TEMPR14[5] ), .D(\R_DATA_TEMPR15[5] ), .Y(OR4_247_Y));
    CFG3 #( .INIT(8'h2) )  CFG3_3 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_3_Y));
    OR4 OR4_518 (.A(\R_DATA_TEMPR44[19] ), .B(\R_DATA_TEMPR45[19] ), 
        .C(\R_DATA_TEMPR46[19] ), .D(\R_DATA_TEMPR47[19] ), .Y(
        OR4_518_Y));
    OR4 OR4_147 (.A(\R_DATA_TEMPR20[5] ), .B(\R_DATA_TEMPR21[5] ), .C(
        \R_DATA_TEMPR22[5] ), .D(\R_DATA_TEMPR23[5] ), .Y(OR4_147_Y));
    OR4 OR4_327 (.A(\R_DATA_TEMPR60[10] ), .B(\R_DATA_TEMPR61[10] ), 
        .C(\R_DATA_TEMPR62[10] ), .D(\R_DATA_TEMPR63[10] ), .Y(
        OR4_327_Y));
    OR4 OR4_120 (.A(\R_DATA_TEMPR16[26] ), .B(\R_DATA_TEMPR17[26] ), 
        .C(\R_DATA_TEMPR18[26] ), .D(\R_DATA_TEMPR19[26] ), .Y(
        OR4_120_Y));
    OR4 OR4_51 (.A(\R_DATA_TEMPR12[34] ), .B(\R_DATA_TEMPR13[34] ), .C(
        \R_DATA_TEMPR14[34] ), .D(\R_DATA_TEMPR15[34] ), .Y(OR4_51_Y));
    CFG1 #( .INIT(2'h1) )  \INVBLKY1[0]  (.A(R_ADDR[10]), .Y(
        \BLKY1[0] ));
    OR4 \OR4_R_DATA[20]  (.A(OR4_585_Y), .B(OR4_774_Y), .C(OR4_331_Y), 
        .D(OR4_28_Y), .Y(R_DATA[20]));
    OR4 OR4_728 (.A(OR4_220_Y), .B(OR4_482_Y), .C(OR4_741_Y), .D(
        OR4_171_Y), .Y(OR4_728_Y));
    OR4 OR4_707 (.A(\R_DATA_TEMPR40[30] ), .B(\R_DATA_TEMPR41[30] ), 
        .C(\R_DATA_TEMPR42[30] ), .D(\R_DATA_TEMPR43[30] ), .Y(
        OR4_707_Y));
    OR4 OR4_704 (.A(\R_DATA_TEMPR40[1] ), .B(\R_DATA_TEMPR41[1] ), .C(
        \R_DATA_TEMPR42[1] ), .D(\R_DATA_TEMPR43[1] ), .Y(OR4_704_Y));
    OR4 OR4_20 (.A(\R_DATA_TEMPR32[1] ), .B(\R_DATA_TEMPR33[1] ), .C(
        \R_DATA_TEMPR34[1] ), .D(\R_DATA_TEMPR35[1] ), .Y(OR4_20_Y));
    OR4 OR4_743 (.A(OR4_478_Y), .B(OR4_668_Y), .C(OR4_122_Y), .D(
        OR4_349_Y), .Y(OR4_743_Y));
    OR4 OR4_777 (.A(\R_DATA_TEMPR60[0] ), .B(\R_DATA_TEMPR61[0] ), .C(
        \R_DATA_TEMPR62[0] ), .D(\R_DATA_TEMPR63[0] ), .Y(OR4_777_Y));
    OR4 OR4_416 (.A(\R_DATA_TEMPR32[22] ), .B(\R_DATA_TEMPR33[22] ), 
        .C(\R_DATA_TEMPR34[22] ), .D(\R_DATA_TEMPR35[22] ), .Y(
        OR4_416_Y));
    OR4 \OR4_R_DATA[26]  (.A(OR4_310_Y), .B(OR4_736_Y), .C(OR4_77_Y), 
        .D(OR4_117_Y), .Y(R_DATA[26]));
    OR4 OR4_774 (.A(OR4_87_Y), .B(OR4_403_Y), .C(OR4_669_Y), .D(
        OR4_368_Y), .Y(OR4_774_Y));
    OR4 OR4_244 (.A(\R_DATA_TEMPR0[3] ), .B(\R_DATA_TEMPR1[3] ), .C(
        \R_DATA_TEMPR2[3] ), .D(\R_DATA_TEMPR3[3] ), .Y(OR4_244_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%12%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R12C0 (
        .A_DOUT({\R_DATA_TEMPR12[39] , \R_DATA_TEMPR12[38] , 
        \R_DATA_TEMPR12[37] , \R_DATA_TEMPR12[36] , 
        \R_DATA_TEMPR12[35] , \R_DATA_TEMPR12[34] , 
        \R_DATA_TEMPR12[33] , \R_DATA_TEMPR12[32] , 
        \R_DATA_TEMPR12[31] , \R_DATA_TEMPR12[30] , 
        \R_DATA_TEMPR12[29] , \R_DATA_TEMPR12[28] , 
        \R_DATA_TEMPR12[27] , \R_DATA_TEMPR12[26] , 
        \R_DATA_TEMPR12[25] , \R_DATA_TEMPR12[24] , 
        \R_DATA_TEMPR12[23] , \R_DATA_TEMPR12[22] , 
        \R_DATA_TEMPR12[21] , \R_DATA_TEMPR12[20] }), .B_DOUT({
        \R_DATA_TEMPR12[19] , \R_DATA_TEMPR12[18] , 
        \R_DATA_TEMPR12[17] , \R_DATA_TEMPR12[16] , 
        \R_DATA_TEMPR12[15] , \R_DATA_TEMPR12[14] , 
        \R_DATA_TEMPR12[13] , \R_DATA_TEMPR12[12] , 
        \R_DATA_TEMPR12[11] , \R_DATA_TEMPR12[10] , 
        \R_DATA_TEMPR12[9] , \R_DATA_TEMPR12[8] , \R_DATA_TEMPR12[7] , 
        \R_DATA_TEMPR12[6] , \R_DATA_TEMPR12[5] , \R_DATA_TEMPR12[4] , 
        \R_DATA_TEMPR12[3] , \R_DATA_TEMPR12[2] , \R_DATA_TEMPR12[1] , 
        \R_DATA_TEMPR12[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_27 (.A(\R_DATA_TEMPR56[18] ), .B(\R_DATA_TEMPR57[18] ), .C(
        \R_DATA_TEMPR58[18] ), .D(\R_DATA_TEMPR59[18] ), .Y(OR4_27_Y));
    OR4 OR4_82 (.A(\R_DATA_TEMPR8[14] ), .B(\R_DATA_TEMPR9[14] ), .C(
        \R_DATA_TEMPR10[14] ), .D(\R_DATA_TEMPR11[14] ), .Y(OR4_82_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R55C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%55%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R55C0 (
        .A_DOUT({\R_DATA_TEMPR55[39] , \R_DATA_TEMPR55[38] , 
        \R_DATA_TEMPR55[37] , \R_DATA_TEMPR55[36] , 
        \R_DATA_TEMPR55[35] , \R_DATA_TEMPR55[34] , 
        \R_DATA_TEMPR55[33] , \R_DATA_TEMPR55[32] , 
        \R_DATA_TEMPR55[31] , \R_DATA_TEMPR55[30] , 
        \R_DATA_TEMPR55[29] , \R_DATA_TEMPR55[28] , 
        \R_DATA_TEMPR55[27] , \R_DATA_TEMPR55[26] , 
        \R_DATA_TEMPR55[25] , \R_DATA_TEMPR55[24] , 
        \R_DATA_TEMPR55[23] , \R_DATA_TEMPR55[22] , 
        \R_DATA_TEMPR55[21] , \R_DATA_TEMPR55[20] }), .B_DOUT({
        \R_DATA_TEMPR55[19] , \R_DATA_TEMPR55[18] , 
        \R_DATA_TEMPR55[17] , \R_DATA_TEMPR55[16] , 
        \R_DATA_TEMPR55[15] , \R_DATA_TEMPR55[14] , 
        \R_DATA_TEMPR55[13] , \R_DATA_TEMPR55[12] , 
        \R_DATA_TEMPR55[11] , \R_DATA_TEMPR55[10] , 
        \R_DATA_TEMPR55[9] , \R_DATA_TEMPR55[8] , \R_DATA_TEMPR55[7] , 
        \R_DATA_TEMPR55[6] , \R_DATA_TEMPR55[5] , \R_DATA_TEMPR55[4] , 
        \R_DATA_TEMPR55[3] , \R_DATA_TEMPR55[2] , \R_DATA_TEMPR55[1] , 
        \R_DATA_TEMPR55[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[55][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[13] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[13] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%30%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R30C0 (
        .A_DOUT({\R_DATA_TEMPR30[39] , \R_DATA_TEMPR30[38] , 
        \R_DATA_TEMPR30[37] , \R_DATA_TEMPR30[36] , 
        \R_DATA_TEMPR30[35] , \R_DATA_TEMPR30[34] , 
        \R_DATA_TEMPR30[33] , \R_DATA_TEMPR30[32] , 
        \R_DATA_TEMPR30[31] , \R_DATA_TEMPR30[30] , 
        \R_DATA_TEMPR30[29] , \R_DATA_TEMPR30[28] , 
        \R_DATA_TEMPR30[27] , \R_DATA_TEMPR30[26] , 
        \R_DATA_TEMPR30[25] , \R_DATA_TEMPR30[24] , 
        \R_DATA_TEMPR30[23] , \R_DATA_TEMPR30[22] , 
        \R_DATA_TEMPR30[21] , \R_DATA_TEMPR30[20] }), .B_DOUT({
        \R_DATA_TEMPR30[19] , \R_DATA_TEMPR30[18] , 
        \R_DATA_TEMPR30[17] , \R_DATA_TEMPR30[16] , 
        \R_DATA_TEMPR30[15] , \R_DATA_TEMPR30[14] , 
        \R_DATA_TEMPR30[13] , \R_DATA_TEMPR30[12] , 
        \R_DATA_TEMPR30[11] , \R_DATA_TEMPR30[10] , 
        \R_DATA_TEMPR30[9] , \R_DATA_TEMPR30[8] , \R_DATA_TEMPR30[7] , 
        \R_DATA_TEMPR30[6] , \R_DATA_TEMPR30[5] , \R_DATA_TEMPR30[4] , 
        \R_DATA_TEMPR30[3] , \R_DATA_TEMPR30[2] , \R_DATA_TEMPR30[1] , 
        \R_DATA_TEMPR30[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[7] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[7] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_128 (.A(\R_DATA_TEMPR40[12] ), .B(\R_DATA_TEMPR41[12] ), 
        .C(\R_DATA_TEMPR42[12] ), .D(\R_DATA_TEMPR43[12] ), .Y(
        OR4_128_Y));
    OR4 OR4_230 (.A(\R_DATA_TEMPR44[18] ), .B(\R_DATA_TEMPR45[18] ), 
        .C(\R_DATA_TEMPR46[18] ), .D(\R_DATA_TEMPR47[18] ), .Y(
        OR4_230_Y));
    OR4 OR4_537 (.A(\R_DATA_TEMPR8[20] ), .B(\R_DATA_TEMPR9[20] ), .C(
        \R_DATA_TEMPR10[20] ), .D(\R_DATA_TEMPR11[20] ), .Y(OR4_537_Y));
    OR4 OR4_182 (.A(\R_DATA_TEMPR28[38] ), .B(\R_DATA_TEMPR29[38] ), 
        .C(\R_DATA_TEMPR30[38] ), .D(\R_DATA_TEMPR31[38] ), .Y(
        OR4_182_Y));
    OR4 OR4_312 (.A(\R_DATA_TEMPR52[33] ), .B(\R_DATA_TEMPR53[33] ), 
        .C(\R_DATA_TEMPR54[33] ), .D(\R_DATA_TEMPR55[33] ), .Y(
        OR4_312_Y));
    OR4 OR4_465 (.A(\R_DATA_TEMPR48[8] ), .B(\R_DATA_TEMPR49[8] ), .C(
        \R_DATA_TEMPR50[8] ), .D(\R_DATA_TEMPR51[8] ), .Y(OR4_465_Y));
    OR4 OR4_551 (.A(\R_DATA_TEMPR60[26] ), .B(\R_DATA_TEMPR61[26] ), 
        .C(\R_DATA_TEMPR62[26] ), .D(\R_DATA_TEMPR63[26] ), .Y(
        OR4_551_Y));
    OR4 OR4_64 (.A(\R_DATA_TEMPR44[8] ), .B(\R_DATA_TEMPR45[8] ), .C(
        \R_DATA_TEMPR46[8] ), .D(\R_DATA_TEMPR47[8] ), .Y(OR4_64_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R39C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%39%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R39C0 (
        .A_DOUT({\R_DATA_TEMPR39[39] , \R_DATA_TEMPR39[38] , 
        \R_DATA_TEMPR39[37] , \R_DATA_TEMPR39[36] , 
        \R_DATA_TEMPR39[35] , \R_DATA_TEMPR39[34] , 
        \R_DATA_TEMPR39[33] , \R_DATA_TEMPR39[32] , 
        \R_DATA_TEMPR39[31] , \R_DATA_TEMPR39[30] , 
        \R_DATA_TEMPR39[29] , \R_DATA_TEMPR39[28] , 
        \R_DATA_TEMPR39[27] , \R_DATA_TEMPR39[26] , 
        \R_DATA_TEMPR39[25] , \R_DATA_TEMPR39[24] , 
        \R_DATA_TEMPR39[23] , \R_DATA_TEMPR39[22] , 
        \R_DATA_TEMPR39[21] , \R_DATA_TEMPR39[20] }), .B_DOUT({
        \R_DATA_TEMPR39[19] , \R_DATA_TEMPR39[18] , 
        \R_DATA_TEMPR39[17] , \R_DATA_TEMPR39[16] , 
        \R_DATA_TEMPR39[15] , \R_DATA_TEMPR39[14] , 
        \R_DATA_TEMPR39[13] , \R_DATA_TEMPR39[12] , 
        \R_DATA_TEMPR39[11] , \R_DATA_TEMPR39[10] , 
        \R_DATA_TEMPR39[9] , \R_DATA_TEMPR39[8] , \R_DATA_TEMPR39[7] , 
        \R_DATA_TEMPR39[6] , \R_DATA_TEMPR39[5] , \R_DATA_TEMPR39[4] , 
        \R_DATA_TEMPR39[3] , \R_DATA_TEMPR39[2] , \R_DATA_TEMPR39[1] , 
        \R_DATA_TEMPR39[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[39][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[9] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[9] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_11 (.A(\R_DATA_TEMPR4[1] ), .B(\R_DATA_TEMPR5[1] ), .C(
        \R_DATA_TEMPR6[1] ), .D(\R_DATA_TEMPR7[1] ), .Y(OR4_11_Y));
    OR4 OR4_639 (.A(\R_DATA_TEMPR52[26] ), .B(\R_DATA_TEMPR53[26] ), 
        .C(\R_DATA_TEMPR54[26] ), .D(\R_DATA_TEMPR55[26] ), .Y(
        OR4_639_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[10]  (.A(CFG3_8_Y), .B(CFG2_3_Y)
        , .Y(\BLKX2[10] ));
    OR4 OR4_345 (.A(\R_DATA_TEMPR28[13] ), .B(\R_DATA_TEMPR29[13] ), 
        .C(\R_DATA_TEMPR30[13] ), .D(\R_DATA_TEMPR31[13] ), .Y(
        OR4_345_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R36C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%36%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R36C0 (
        .A_DOUT({\R_DATA_TEMPR36[39] , \R_DATA_TEMPR36[38] , 
        \R_DATA_TEMPR36[37] , \R_DATA_TEMPR36[36] , 
        \R_DATA_TEMPR36[35] , \R_DATA_TEMPR36[34] , 
        \R_DATA_TEMPR36[33] , \R_DATA_TEMPR36[32] , 
        \R_DATA_TEMPR36[31] , \R_DATA_TEMPR36[30] , 
        \R_DATA_TEMPR36[29] , \R_DATA_TEMPR36[28] , 
        \R_DATA_TEMPR36[27] , \R_DATA_TEMPR36[26] , 
        \R_DATA_TEMPR36[25] , \R_DATA_TEMPR36[24] , 
        \R_DATA_TEMPR36[23] , \R_DATA_TEMPR36[22] , 
        \R_DATA_TEMPR36[21] , \R_DATA_TEMPR36[20] }), .B_DOUT({
        \R_DATA_TEMPR36[19] , \R_DATA_TEMPR36[18] , 
        \R_DATA_TEMPR36[17] , \R_DATA_TEMPR36[16] , 
        \R_DATA_TEMPR36[15] , \R_DATA_TEMPR36[14] , 
        \R_DATA_TEMPR36[13] , \R_DATA_TEMPR36[12] , 
        \R_DATA_TEMPR36[11] , \R_DATA_TEMPR36[10] , 
        \R_DATA_TEMPR36[9] , \R_DATA_TEMPR36[8] , \R_DATA_TEMPR36[7] , 
        \R_DATA_TEMPR36[6] , \R_DATA_TEMPR36[5] , \R_DATA_TEMPR36[4] , 
        \R_DATA_TEMPR36[3] , \R_DATA_TEMPR36[2] , \R_DATA_TEMPR36[1] , 
        \R_DATA_TEMPR36[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[36][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[9] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[9] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_236 (.A(\R_DATA_TEMPR48[37] ), .B(\R_DATA_TEMPR49[37] ), 
        .C(\R_DATA_TEMPR50[37] ), .D(\R_DATA_TEMPR51[37] ), .Y(
        OR4_236_Y));
    OR4 OR4_73 (.A(OR4_430_Y), .B(OR4_544_Y), .C(OR4_535_Y), .D(
        OR4_104_Y), .Y(OR4_73_Y));
    OR4 OR4_195 (.A(\R_DATA_TEMPR8[6] ), .B(\R_DATA_TEMPR9[6] ), .C(
        \R_DATA_TEMPR10[6] ), .D(\R_DATA_TEMPR11[6] ), .Y(OR4_195_Y));
    OR4 OR4_252 (.A(\R_DATA_TEMPR20[30] ), .B(\R_DATA_TEMPR21[30] ), 
        .C(\R_DATA_TEMPR22[30] ), .D(\R_DATA_TEMPR23[30] ), .Y(
        OR4_252_Y));
    OR4 OR4_289 (.A(\R_DATA_TEMPR40[22] ), .B(\R_DATA_TEMPR41[22] ), 
        .C(\R_DATA_TEMPR42[22] ), .D(\R_DATA_TEMPR43[22] ), .Y(
        OR4_289_Y));
    OR4 OR4_497 (.A(\R_DATA_TEMPR24[23] ), .B(\R_DATA_TEMPR25[23] ), 
        .C(\R_DATA_TEMPR26[23] ), .D(\R_DATA_TEMPR27[23] ), .Y(
        OR4_497_Y));
    OR4 OR4_634 (.A(\R_DATA_TEMPR28[5] ), .B(\R_DATA_TEMPR29[5] ), .C(
        \R_DATA_TEMPR30[5] ), .D(\R_DATA_TEMPR31[5] ), .Y(OR4_634_Y));
    OR4 OR4_464 (.A(\R_DATA_TEMPR40[28] ), .B(\R_DATA_TEMPR41[28] ), 
        .C(\R_DATA_TEMPR42[28] ), .D(\R_DATA_TEMPR43[28] ), .Y(
        OR4_464_Y));
    OR4 OR4_210 (.A(OR4_685_Y), .B(OR4_601_Y), .C(OR4_307_Y), .D(
        OR4_558_Y), .Y(OR4_210_Y));
    OR4 OR4_742 (.A(\R_DATA_TEMPR52[23] ), .B(\R_DATA_TEMPR53[23] ), 
        .C(\R_DATA_TEMPR54[23] ), .D(\R_DATA_TEMPR55[23] ), .Y(
        OR4_742_Y));
    OR4 OR4_517 (.A(\R_DATA_TEMPR8[23] ), .B(\R_DATA_TEMPR9[23] ), .C(
        \R_DATA_TEMPR10[23] ), .D(\R_DATA_TEMPR11[23] ), .Y(OR4_517_Y));
    OR4 OR4_350 (.A(\R_DATA_TEMPR48[28] ), .B(\R_DATA_TEMPR49[28] ), 
        .C(\R_DATA_TEMPR50[28] ), .D(\R_DATA_TEMPR51[28] ), .Y(
        OR4_350_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[1]  (.A(CFG3_4_Y), .B(CFG2_2_Y), 
        .Y(\BLKX2[1] ));
    OR4 OR4_366 (.A(\R_DATA_TEMPR32[3] ), .B(\R_DATA_TEMPR33[3] ), .C(
        \R_DATA_TEMPR34[3] ), .D(\R_DATA_TEMPR35[3] ), .Y(OR4_366_Y));
    OR4 OR4_295 (.A(\R_DATA_TEMPR36[27] ), .B(\R_DATA_TEMPR37[27] ), 
        .C(\R_DATA_TEMPR38[27] ), .D(\R_DATA_TEMPR39[27] ), .Y(
        OR4_295_Y));
    OR4 OR4_645 (.A(\R_DATA_TEMPR48[29] ), .B(\R_DATA_TEMPR49[29] ), 
        .C(\R_DATA_TEMPR50[29] ), .D(\R_DATA_TEMPR51[29] ), .Y(
        OR4_645_Y));
    OR4 OR4_619 (.A(\R_DATA_TEMPR32[2] ), .B(\R_DATA_TEMPR33[2] ), .C(
        \R_DATA_TEMPR34[2] ), .D(\R_DATA_TEMPR35[2] ), .Y(OR4_619_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[13]  (.A(CFG3_14_Y), .B(
        CFG2_3_Y), .Y(\BLKX2[13] ));
    OR4 OR4_35 (.A(\R_DATA_TEMPR52[22] ), .B(\R_DATA_TEMPR53[22] ), .C(
        \R_DATA_TEMPR54[22] ), .D(\R_DATA_TEMPR55[22] ), .Y(OR4_35_Y));
    OR4 OR4_405 (.A(\R_DATA_TEMPR60[28] ), .B(\R_DATA_TEMPR61[28] ), 
        .C(\R_DATA_TEMPR62[28] ), .D(\R_DATA_TEMPR63[28] ), .Y(
        OR4_405_Y));
    OR4 OR4_216 (.A(OR4_700_Y), .B(OR4_445_Y), .C(OR4_708_Y), .D(
        OR4_412_Y), .Y(OR4_216_Y));
    OR4 OR4_71 (.A(\R_DATA_TEMPR36[24] ), .B(\R_DATA_TEMPR37[24] ), .C(
        \R_DATA_TEMPR38[24] ), .D(\R_DATA_TEMPR39[24] ), .Y(OR4_71_Y));
    OR4 OR4_475 (.A(\R_DATA_TEMPR44[37] ), .B(\R_DATA_TEMPR45[37] ), 
        .C(\R_DATA_TEMPR46[37] ), .D(\R_DATA_TEMPR47[37] ), .Y(
        OR4_475_Y));
    OR4 OR4_125 (.A(\R_DATA_TEMPR56[1] ), .B(\R_DATA_TEMPR57[1] ), .C(
        \R_DATA_TEMPR58[1] ), .D(\R_DATA_TEMPR59[1] ), .Y(OR4_125_Y));
    OR4 OR4_493 (.A(\R_DATA_TEMPR12[7] ), .B(\R_DATA_TEMPR13[7] ), .C(
        \R_DATA_TEMPR14[7] ), .D(\R_DATA_TEMPR15[7] ), .Y(OR4_493_Y));
    OR4 OR4_691 (.A(\R_DATA_TEMPR0[26] ), .B(\R_DATA_TEMPR1[26] ), .C(
        \R_DATA_TEMPR2[26] ), .D(\R_DATA_TEMPR3[26] ), .Y(OR4_691_Y));
    OR4 OR4_614 (.A(\R_DATA_TEMPR40[19] ), .B(\R_DATA_TEMPR41[19] ), 
        .C(\R_DATA_TEMPR42[19] ), .D(\R_DATA_TEMPR43[19] ), .Y(
        OR4_614_Y));
    OR4 OR4_427 (.A(\R_DATA_TEMPR56[32] ), .B(\R_DATA_TEMPR57[32] ), 
        .C(\R_DATA_TEMPR58[32] ), .D(\R_DATA_TEMPR59[32] ), .Y(
        OR4_427_Y));
    OR4 OR4_787 (.A(\R_DATA_TEMPR20[13] ), .B(\R_DATA_TEMPR21[13] ), 
        .C(\R_DATA_TEMPR22[13] ), .D(\R_DATA_TEMPR23[13] ), .Y(
        OR4_787_Y));
    OR4 OR4_298 (.A(OR4_47_Y), .B(OR4_202_Y), .C(OR4_319_Y), .D(
        OR4_230_Y), .Y(OR4_298_Y));
    OR4 \OR4_R_DATA[27]  (.A(OR4_100_Y), .B(OR4_483_Y), .C(OR4_689_Y), 
        .D(OR4_768_Y), .Y(R_DATA[27]));
    OR4 OR4_784 (.A(\R_DATA_TEMPR4[29] ), .B(\R_DATA_TEMPR5[29] ), .C(
        \R_DATA_TEMPR6[29] ), .D(\R_DATA_TEMPR7[29] ), .Y(OR4_784_Y));
    OR4 OR4_28 (.A(OR4_250_Y), .B(OR4_106_Y), .C(OR4_782_Y), .D(
        OR4_580_Y), .Y(OR4_28_Y));
    OR4 OR4_640 (.A(\R_DATA_TEMPR4[5] ), .B(\R_DATA_TEMPR5[5] ), .C(
        \R_DATA_TEMPR6[5] ), .D(\R_DATA_TEMPR7[5] ), .Y(OR4_640_Y));
    OR4 OR4_164 (.A(\R_DATA_TEMPR40[9] ), .B(\R_DATA_TEMPR41[9] ), .C(
        \R_DATA_TEMPR42[9] ), .D(\R_DATA_TEMPR43[9] ), .Y(OR4_164_Y));
    OR4 OR4_404 (.A(\R_DATA_TEMPR8[38] ), .B(\R_DATA_TEMPR9[38] ), .C(
        \R_DATA_TEMPR10[38] ), .D(\R_DATA_TEMPR11[38] ), .Y(OR4_404_Y));
    OR4 OR4_225 (.A(\R_DATA_TEMPR12[2] ), .B(\R_DATA_TEMPR13[2] ), .C(
        \R_DATA_TEMPR14[2] ), .D(\R_DATA_TEMPR15[2] ), .Y(OR4_225_Y));
    CFG2 #( .INIT(4'h2) )  CFG2_2 (.A(W_EN), .B(W_ADDR[14]), .Y(
        CFG2_2_Y));
    OR4 OR4_555 (.A(\R_DATA_TEMPR48[27] ), .B(\R_DATA_TEMPR49[27] ), 
        .C(\R_DATA_TEMPR50[27] ), .D(\R_DATA_TEMPR51[27] ), .Y(
        OR4_555_Y));
    OR4 OR4_347 (.A(\R_DATA_TEMPR48[24] ), .B(\R_DATA_TEMPR49[24] ), 
        .C(\R_DATA_TEMPR50[24] ), .D(\R_DATA_TEMPR51[24] ), .Y(
        OR4_347_Y));
    OR4 OR4_140 (.A(\R_DATA_TEMPR56[0] ), .B(\R_DATA_TEMPR57[0] ), .C(
        \R_DATA_TEMPR58[0] ), .D(\R_DATA_TEMPR59[0] ), .Y(OR4_140_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R62C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%62%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R62C0 (
        .A_DOUT({\R_DATA_TEMPR62[39] , \R_DATA_TEMPR62[38] , 
        \R_DATA_TEMPR62[37] , \R_DATA_TEMPR62[36] , 
        \R_DATA_TEMPR62[35] , \R_DATA_TEMPR62[34] , 
        \R_DATA_TEMPR62[33] , \R_DATA_TEMPR62[32] , 
        \R_DATA_TEMPR62[31] , \R_DATA_TEMPR62[30] , 
        \R_DATA_TEMPR62[29] , \R_DATA_TEMPR62[28] , 
        \R_DATA_TEMPR62[27] , \R_DATA_TEMPR62[26] , 
        \R_DATA_TEMPR62[25] , \R_DATA_TEMPR62[24] , 
        \R_DATA_TEMPR62[23] , \R_DATA_TEMPR62[22] , 
        \R_DATA_TEMPR62[21] , \R_DATA_TEMPR62[20] }), .B_DOUT({
        \R_DATA_TEMPR62[19] , \R_DATA_TEMPR62[18] , 
        \R_DATA_TEMPR62[17] , \R_DATA_TEMPR62[16] , 
        \R_DATA_TEMPR62[15] , \R_DATA_TEMPR62[14] , 
        \R_DATA_TEMPR62[13] , \R_DATA_TEMPR62[12] , 
        \R_DATA_TEMPR62[11] , \R_DATA_TEMPR62[10] , 
        \R_DATA_TEMPR62[9] , \R_DATA_TEMPR62[8] , \R_DATA_TEMPR62[7] , 
        \R_DATA_TEMPR62[6] , \R_DATA_TEMPR62[5] , \R_DATA_TEMPR62[4] , 
        \R_DATA_TEMPR62[3] , \R_DATA_TEMPR62[2] , \R_DATA_TEMPR62[1] , 
        \R_DATA_TEMPR62[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[62][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[15] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[15] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_474 (.A(\R_DATA_TEMPR56[3] ), .B(\R_DATA_TEMPR57[3] ), .C(
        \R_DATA_TEMPR58[3] ), .D(\R_DATA_TEMPR59[3] ), .Y(OR4_474_Y));
    OR4 OR4_306 (.A(\R_DATA_TEMPR60[22] ), .B(\R_DATA_TEMPR61[22] ), 
        .C(\R_DATA_TEMPR62[22] ), .D(\R_DATA_TEMPR63[22] ), .Y(
        OR4_306_Y));
    OR4 OR4_748 (.A(\R_DATA_TEMPR0[13] ), .B(\R_DATA_TEMPR1[13] ), .C(
        \R_DATA_TEMPR2[13] ), .D(\R_DATA_TEMPR3[13] ), .Y(OR4_748_Y));
    OR4 OR4_653 (.A(\R_DATA_TEMPR24[16] ), .B(\R_DATA_TEMPR25[16] ), 
        .C(\R_DATA_TEMPR26[16] ), .D(\R_DATA_TEMPR27[16] ), .Y(
        OR4_653_Y));
    CFG2 #( .INIT(4'h8) )  CFG2_3 (.A(W_EN), .B(W_ADDR[14]), .Y(
        CFG2_3_Y));
    OR4 OR4_376 (.A(\R_DATA_TEMPR52[16] ), .B(\R_DATA_TEMPR53[16] ), 
        .C(\R_DATA_TEMPR54[16] ), .D(\R_DATA_TEMPR55[16] ), .Y(
        OR4_376_Y));
    OR4 OR4_761 (.A(\R_DATA_TEMPR52[14] ), .B(\R_DATA_TEMPR53[14] ), 
        .C(\R_DATA_TEMPR54[14] ), .D(\R_DATA_TEMPR55[14] ), .Y(
        OR4_761_Y));
    OR4 OR4_423 (.A(OR4_41_Y), .B(OR4_761_Y), .C(OR4_23_Y), .D(
        OR4_775_Y), .Y(OR4_423_Y));
    OR4 OR4_621 (.A(\R_DATA_TEMPR28[14] ), .B(\R_DATA_TEMPR29[14] ), 
        .C(\R_DATA_TEMPR30[14] ), .D(\R_DATA_TEMPR31[14] ), .Y(
        OR4_621_Y));
    OR4 OR4_84 (.A(\R_DATA_TEMPR32[11] ), .B(\R_DATA_TEMPR33[11] ), .C(
        \R_DATA_TEMPR34[11] ), .D(\R_DATA_TEMPR35[11] ), .Y(OR4_84_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[13]  (.A(CFG3_6_Y), .B(CFG2_1_Y)
        , .Y(\BLKY2[13] ));
    OR4 OR4_148 (.A(\R_DATA_TEMPR16[22] ), .B(\R_DATA_TEMPR17[22] ), 
        .C(\R_DATA_TEMPR18[22] ), .D(\R_DATA_TEMPR19[22] ), .Y(
        OR4_148_Y));
    OR4 OR4_228 (.A(\R_DATA_TEMPR44[14] ), .B(\R_DATA_TEMPR45[14] ), 
        .C(\R_DATA_TEMPR46[14] ), .D(\R_DATA_TEMPR47[14] ), .Y(
        OR4_228_Y));
    OR4 OR4_566 (.A(\R_DATA_TEMPR8[5] ), .B(\R_DATA_TEMPR9[5] ), .C(
        \R_DATA_TEMPR10[5] ), .D(\R_DATA_TEMPR11[5] ), .Y(OR4_566_Y));
    OR4 OR4_591 (.A(\R_DATA_TEMPR44[28] ), .B(\R_DATA_TEMPR45[28] ), 
        .C(\R_DATA_TEMPR46[28] ), .D(\R_DATA_TEMPR47[28] ), .Y(
        OR4_591_Y));
    CFG3 #( .INIT(8'h10) )  CFG3_4 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_4_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[9]  (.A(CFG3_4_Y), .B(CFG2_3_Y), 
        .Y(\BLKX2[9] ));
    OR4 OR4_153 (.A(\R_DATA_TEMPR16[10] ), .B(\R_DATA_TEMPR17[10] ), 
        .C(\R_DATA_TEMPR18[10] ), .D(\R_DATA_TEMPR19[10] ), .Y(
        OR4_153_Y));
    OR4 OR4_9 (.A(OR4_361_Y), .B(OR4_797_Y), .C(OR4_274_Y), .D(
        OR4_773_Y), .Y(OR4_9_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%27%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R27C0 (
        .A_DOUT({\R_DATA_TEMPR27[39] , \R_DATA_TEMPR27[38] , 
        \R_DATA_TEMPR27[37] , \R_DATA_TEMPR27[36] , 
        \R_DATA_TEMPR27[35] , \R_DATA_TEMPR27[34] , 
        \R_DATA_TEMPR27[33] , \R_DATA_TEMPR27[32] , 
        \R_DATA_TEMPR27[31] , \R_DATA_TEMPR27[30] , 
        \R_DATA_TEMPR27[29] , \R_DATA_TEMPR27[28] , 
        \R_DATA_TEMPR27[27] , \R_DATA_TEMPR27[26] , 
        \R_DATA_TEMPR27[25] , \R_DATA_TEMPR27[24] , 
        \R_DATA_TEMPR27[23] , \R_DATA_TEMPR27[22] , 
        \R_DATA_TEMPR27[21] , \R_DATA_TEMPR27[20] }), .B_DOUT({
        \R_DATA_TEMPR27[19] , \R_DATA_TEMPR27[18] , 
        \R_DATA_TEMPR27[17] , \R_DATA_TEMPR27[16] , 
        \R_DATA_TEMPR27[15] , \R_DATA_TEMPR27[14] , 
        \R_DATA_TEMPR27[13] , \R_DATA_TEMPR27[12] , 
        \R_DATA_TEMPR27[11] , \R_DATA_TEMPR27[10] , 
        \R_DATA_TEMPR27[9] , \R_DATA_TEMPR27[8] , \R_DATA_TEMPR27[7] , 
        \R_DATA_TEMPR27[6] , \R_DATA_TEMPR27[5] , \R_DATA_TEMPR27[4] , 
        \R_DATA_TEMPR27[3] , \R_DATA_TEMPR27[2] , \R_DATA_TEMPR27[1] , 
        \R_DATA_TEMPR27[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[6] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[6] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_231 (.A(OR4_568_Y), .B(OR4_486_Y), .C(OR4_550_Y), .D(
        OR4_564_Y), .Y(OR4_231_Y));
    OR4 OR4_104 (.A(\R_DATA_TEMPR28[19] ), .B(\R_DATA_TEMPR29[19] ), 
        .C(\R_DATA_TEMPR30[19] ), .D(\R_DATA_TEMPR31[19] ), .Y(
        OR4_104_Y));
    OR4 OR4_292 (.A(\R_DATA_TEMPR4[28] ), .B(\R_DATA_TEMPR5[28] ), .C(
        \R_DATA_TEMPR6[28] ), .D(\R_DATA_TEMPR7[28] ), .Y(OR4_292_Y));
    CFG3 #( .INIT(8'h8) )  CFG3_5 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_5_Y));
    OR4 OR4_174 (.A(\R_DATA_TEMPR12[9] ), .B(\R_DATA_TEMPR13[9] ), .C(
        \R_DATA_TEMPR14[9] ), .D(\R_DATA_TEMPR15[9] ), .Y(OR4_174_Y));
    OR4 OR4_485 (.A(OR4_148_Y), .B(OR4_326_Y), .C(OR4_588_Y), .D(
        OR4_300_Y), .Y(OR4_485_Y));
    OR4 OR4_568 (.A(\R_DATA_TEMPR48[13] ), .B(\R_DATA_TEMPR49[13] ), 
        .C(\R_DATA_TEMPR50[13] ), .D(\R_DATA_TEMPR51[13] ), .Y(
        OR4_568_Y));
    OR4 OR4_532 (.A(\R_DATA_TEMPR16[8] ), .B(\R_DATA_TEMPR17[8] ), .C(
        \R_DATA_TEMPR18[8] ), .D(\R_DATA_TEMPR19[8] ), .Y(OR4_532_Y));
    OR4 OR4_56 (.A(\R_DATA_TEMPR56[11] ), .B(\R_DATA_TEMPR57[11] ), .C(
        \R_DATA_TEMPR58[11] ), .D(\R_DATA_TEMPR59[11] ), .Y(OR4_56_Y));
    OR4 OR4_390 (.A(\R_DATA_TEMPR20[31] ), .B(\R_DATA_TEMPR21[31] ), 
        .C(\R_DATA_TEMPR22[31] ), .D(\R_DATA_TEMPR23[31] ), .Y(
        OR4_390_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%15%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R15C0 (
        .A_DOUT({\R_DATA_TEMPR15[39] , \R_DATA_TEMPR15[38] , 
        \R_DATA_TEMPR15[37] , \R_DATA_TEMPR15[36] , 
        \R_DATA_TEMPR15[35] , \R_DATA_TEMPR15[34] , 
        \R_DATA_TEMPR15[33] , \R_DATA_TEMPR15[32] , 
        \R_DATA_TEMPR15[31] , \R_DATA_TEMPR15[30] , 
        \R_DATA_TEMPR15[29] , \R_DATA_TEMPR15[28] , 
        \R_DATA_TEMPR15[27] , \R_DATA_TEMPR15[26] , 
        \R_DATA_TEMPR15[25] , \R_DATA_TEMPR15[24] , 
        \R_DATA_TEMPR15[23] , \R_DATA_TEMPR15[22] , 
        \R_DATA_TEMPR15[21] , \R_DATA_TEMPR15[20] }), .B_DOUT({
        \R_DATA_TEMPR15[19] , \R_DATA_TEMPR15[18] , 
        \R_DATA_TEMPR15[17] , \R_DATA_TEMPR15[16] , 
        \R_DATA_TEMPR15[15] , \R_DATA_TEMPR15[14] , 
        \R_DATA_TEMPR15[13] , \R_DATA_TEMPR15[12] , 
        \R_DATA_TEMPR15[11] , \R_DATA_TEMPR15[10] , 
        \R_DATA_TEMPR15[9] , \R_DATA_TEMPR15[8] , \R_DATA_TEMPR15[7] , 
        \R_DATA_TEMPR15[6] , \R_DATA_TEMPR15[5] , \R_DATA_TEMPR15[4] , 
        \R_DATA_TEMPR15[3] , \R_DATA_TEMPR15[2] , \R_DATA_TEMPR15[1] , 
        \R_DATA_TEMPR15[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_701 (.A(\R_DATA_TEMPR0[38] ), .B(\R_DATA_TEMPR1[38] ), .C(
        \R_DATA_TEMPR2[38] ), .D(\R_DATA_TEMPR3[38] ), .Y(OR4_701_Y));
    OR4 \OR4_R_DATA[2]  (.A(OR4_441_Y), .B(OR4_397_Y), .C(OR4_549_Y), 
        .D(OR4_610_Y), .Y(R_DATA[2]));
    OR4 OR4_521 (.A(\R_DATA_TEMPR28[21] ), .B(\R_DATA_TEMPR29[21] ), 
        .C(\R_DATA_TEMPR30[21] ), .D(\R_DATA_TEMPR31[21] ), .Y(
        OR4_521_Y));
    OR4 OR4_771 (.A(\R_DATA_TEMPR16[15] ), .B(\R_DATA_TEMPR17[15] ), 
        .C(\R_DATA_TEMPR18[15] ), .D(\R_DATA_TEMPR19[15] ), .Y(
        OR4_771_Y));
    OR4 OR4_152 (.A(OR4_54_Y), .B(OR4_632_Y), .C(OR4_89_Y), .D(
        OR4_314_Y), .Y(OR4_152_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R32C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%32%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R32C0 (
        .A_DOUT({\R_DATA_TEMPR32[39] , \R_DATA_TEMPR32[38] , 
        \R_DATA_TEMPR32[37] , \R_DATA_TEMPR32[36] , 
        \R_DATA_TEMPR32[35] , \R_DATA_TEMPR32[34] , 
        \R_DATA_TEMPR32[33] , \R_DATA_TEMPR32[32] , 
        \R_DATA_TEMPR32[31] , \R_DATA_TEMPR32[30] , 
        \R_DATA_TEMPR32[29] , \R_DATA_TEMPR32[28] , 
        \R_DATA_TEMPR32[27] , \R_DATA_TEMPR32[26] , 
        \R_DATA_TEMPR32[25] , \R_DATA_TEMPR32[24] , 
        \R_DATA_TEMPR32[23] , \R_DATA_TEMPR32[22] , 
        \R_DATA_TEMPR32[21] , \R_DATA_TEMPR32[20] }), .B_DOUT({
        \R_DATA_TEMPR32[19] , \R_DATA_TEMPR32[18] , 
        \R_DATA_TEMPR32[17] , \R_DATA_TEMPR32[16] , 
        \R_DATA_TEMPR32[15] , \R_DATA_TEMPR32[14] , 
        \R_DATA_TEMPR32[13] , \R_DATA_TEMPR32[12] , 
        \R_DATA_TEMPR32[11] , \R_DATA_TEMPR32[10] , 
        \R_DATA_TEMPR32[9] , \R_DATA_TEMPR32[8] , \R_DATA_TEMPR32[7] , 
        \R_DATA_TEMPR32[6] , \R_DATA_TEMPR32[5] , \R_DATA_TEMPR32[4] , 
        \R_DATA_TEMPR32[3] , \R_DATA_TEMPR32[2] , \R_DATA_TEMPR32[1] , 
        \R_DATA_TEMPR32[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[32][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[8] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[8] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_466 (.A(\R_DATA_TEMPR24[6] ), .B(\R_DATA_TEMPR25[6] ), .C(
        \R_DATA_TEMPR26[6] ), .D(\R_DATA_TEMPR27[6] ), .Y(OR4_466_Y));
    OR4 OR4_39 (.A(\R_DATA_TEMPR44[12] ), .B(\R_DATA_TEMPR45[12] ), .C(
        \R_DATA_TEMPR46[12] ), .D(\R_DATA_TEMPR47[12] ), .Y(OR4_39_Y));
    OR4 OR4_534 (.A(OR4_81_Y), .B(OR4_3_Y), .C(OR4_56_Y), .D(OR4_263_Y)
        , .Y(OR4_534_Y));
    OR4 OR4_506 (.A(\R_DATA_TEMPR60[21] ), .B(\R_DATA_TEMPR61[21] ), 
        .C(\R_DATA_TEMPR62[21] ), .D(\R_DATA_TEMPR63[21] ), .Y(
        OR4_506_Y));
    OR4 OR4_211 (.A(\R_DATA_TEMPR32[26] ), .B(\R_DATA_TEMPR33[26] ), 
        .C(\R_DATA_TEMPR34[26] ), .D(\R_DATA_TEMPR35[26] ), .Y(
        OR4_211_Y));
    OR4 OR4_484 (.A(OR4_748_Y), .B(OR4_595_Y), .C(OR4_578_Y), .D(
        OR4_281_Y), .Y(OR4_484_Y));
    OR4 OR4_576 (.A(\R_DATA_TEMPR4[32] ), .B(\R_DATA_TEMPR5[32] ), .C(
        \R_DATA_TEMPR6[32] ), .D(\R_DATA_TEMPR7[32] ), .Y(OR4_576_Y));
    OR4 OR4_145 (.A(\R_DATA_TEMPR60[32] ), .B(\R_DATA_TEMPR61[32] ), 
        .C(\R_DATA_TEMPR62[32] ), .D(\R_DATA_TEMPR63[32] ), .Y(
        OR4_145_Y));
    OR4 OR4_362 (.A(\R_DATA_TEMPR32[6] ), .B(\R_DATA_TEMPR33[6] ), .C(
        \R_DATA_TEMPR34[6] ), .D(\R_DATA_TEMPR35[6] ), .Y(OR4_362_Y));
    OR4 OR4_222 (.A(\R_DATA_TEMPR8[18] ), .B(\R_DATA_TEMPR9[18] ), .C(
        \R_DATA_TEMPR10[18] ), .D(\R_DATA_TEMPR11[18] ), .Y(OR4_222_Y));
    OR4 OR4_16 (.A(\R_DATA_TEMPR36[12] ), .B(\R_DATA_TEMPR37[12] ), .C(
        \R_DATA_TEMPR38[12] ), .D(\R_DATA_TEMPR39[12] ), .Y(OR4_16_Y));
    OR4 OR4_386 (.A(\R_DATA_TEMPR56[9] ), .B(\R_DATA_TEMPR57[9] ), .C(
        \R_DATA_TEMPR58[9] ), .D(\R_DATA_TEMPR59[9] ), .Y(OR4_386_Y));
    OR4 OR4_447 (.A(\R_DATA_TEMPR8[9] ), .B(\R_DATA_TEMPR9[9] ), .C(
        \R_DATA_TEMPR10[9] ), .D(\R_DATA_TEMPR11[9] ), .Y(OR4_447_Y));
    OR4 OR4_259 (.A(\R_DATA_TEMPR0[9] ), .B(\R_DATA_TEMPR1[9] ), .C(
        \R_DATA_TEMPR2[9] ), .D(\R_DATA_TEMPR3[9] ), .Y(OR4_259_Y));
    OR4 OR4_4 (.A(\R_DATA_TEMPR32[36] ), .B(\R_DATA_TEMPR33[36] ), .C(
        \R_DATA_TEMPR34[36] ), .D(\R_DATA_TEMPR35[36] ), .Y(OR4_4_Y));
    OR4 OR4_331 (.A(OR4_487_Y), .B(OR4_780_Y), .C(OR4_359_Y), .D(
        OR4_481_Y), .Y(OR4_331_Y));
    OR4 OR4_512 (.A(OR4_658_Y), .B(OR4_330_Y), .C(OR4_494_Y), .D(
        OR4_93_Y), .Y(OR4_512_Y));
    OR4 OR4_320 (.A(\R_DATA_TEMPR44[23] ), .B(\R_DATA_TEMPR45[23] ), 
        .C(\R_DATA_TEMPR46[23] ), .D(\R_DATA_TEMPR47[23] ), .Y(
        OR4_320_Y));
    OR4 OR4_430 (.A(\R_DATA_TEMPR16[19] ), .B(\R_DATA_TEMPR17[19] ), 
        .C(\R_DATA_TEMPR18[19] ), .D(\R_DATA_TEMPR19[19] ), .Y(
        OR4_430_Y));
    OR4 \OR4_R_DATA[14]  (.A(OR4_757_Y), .B(OR4_480_Y), .C(OR4_62_Y), 
        .D(OR4_423_Y), .Y(R_DATA[14]));
    OR4 OR4_595 (.A(\R_DATA_TEMPR4[13] ), .B(\R_DATA_TEMPR5[13] ), .C(
        \R_DATA_TEMPR6[13] ), .D(\R_DATA_TEMPR7[13] ), .Y(OR4_595_Y));
    OR4 OR4_245 (.A(\R_DATA_TEMPR4[4] ), .B(\R_DATA_TEMPR5[4] ), .C(
        \R_DATA_TEMPR6[4] ), .D(\R_DATA_TEMPR7[4] ), .Y(OR4_245_Y));
    OR4 OR4_508 (.A(\R_DATA_TEMPR0[29] ), .B(\R_DATA_TEMPR1[29] ), .C(
        \R_DATA_TEMPR2[29] ), .D(\R_DATA_TEMPR3[29] ), .Y(OR4_508_Y));
    OR4 OR4_50 (.A(\R_DATA_TEMPR40[31] ), .B(\R_DATA_TEMPR41[31] ), .C(
        \R_DATA_TEMPR42[31] ), .D(\R_DATA_TEMPR43[31] ), .Y(OR4_50_Y));
    OR4 OR4_514 (.A(\R_DATA_TEMPR28[10] ), .B(\R_DATA_TEMPR29[10] ), 
        .C(\R_DATA_TEMPR30[10] ), .D(\R_DATA_TEMPR31[10] ), .Y(
        OR4_514_Y));
    OR4 OR4_578 (.A(\R_DATA_TEMPR8[13] ), .B(\R_DATA_TEMPR9[13] ), .C(
        \R_DATA_TEMPR10[13] ), .D(\R_DATA_TEMPR11[13] ), .Y(OR4_578_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R57C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%57%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R57C0 (
        .A_DOUT({\R_DATA_TEMPR57[39] , \R_DATA_TEMPR57[38] , 
        \R_DATA_TEMPR57[37] , \R_DATA_TEMPR57[36] , 
        \R_DATA_TEMPR57[35] , \R_DATA_TEMPR57[34] , 
        \R_DATA_TEMPR57[33] , \R_DATA_TEMPR57[32] , 
        \R_DATA_TEMPR57[31] , \R_DATA_TEMPR57[30] , 
        \R_DATA_TEMPR57[29] , \R_DATA_TEMPR57[28] , 
        \R_DATA_TEMPR57[27] , \R_DATA_TEMPR57[26] , 
        \R_DATA_TEMPR57[25] , \R_DATA_TEMPR57[24] , 
        \R_DATA_TEMPR57[23] , \R_DATA_TEMPR57[22] , 
        \R_DATA_TEMPR57[21] , \R_DATA_TEMPR57[20] }), .B_DOUT({
        \R_DATA_TEMPR57[19] , \R_DATA_TEMPR57[18] , 
        \R_DATA_TEMPR57[17] , \R_DATA_TEMPR57[16] , 
        \R_DATA_TEMPR57[15] , \R_DATA_TEMPR57[14] , 
        \R_DATA_TEMPR57[13] , \R_DATA_TEMPR57[12] , 
        \R_DATA_TEMPR57[11] , \R_DATA_TEMPR57[10] , 
        \R_DATA_TEMPR57[9] , \R_DATA_TEMPR57[8] , \R_DATA_TEMPR57[7] , 
        \R_DATA_TEMPR57[6] , \R_DATA_TEMPR57[5] , \R_DATA_TEMPR57[4] , 
        \R_DATA_TEMPR57[3] , \R_DATA_TEMPR57[2] , \R_DATA_TEMPR57[1] , 
        \R_DATA_TEMPR57[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[57][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[14] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[14] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_693 (.A(\R_DATA_TEMPR16[14] ), .B(\R_DATA_TEMPR17[14] ), 
        .C(\R_DATA_TEMPR18[14] ), .D(\R_DATA_TEMPR19[14] ), .Y(
        OR4_693_Y));
    OR4 OR4_57 (.A(\R_DATA_TEMPR24[33] ), .B(\R_DATA_TEMPR25[33] ), .C(
        \R_DATA_TEMPR26[33] ), .D(\R_DATA_TEMPR27[33] ), .Y(OR4_57_Y));
    OR4 OR4_32 (.A(\R_DATA_TEMPR36[33] ), .B(\R_DATA_TEMPR37[33] ), .C(
        \R_DATA_TEMPR38[33] ), .D(\R_DATA_TEMPR39[33] ), .Y(OR4_32_Y));
    OR4 OR4_260 (.A(\R_DATA_TEMPR48[17] ), .B(\R_DATA_TEMPR49[17] ), 
        .C(\R_DATA_TEMPR50[17] ), .D(\R_DATA_TEMPR51[17] ), .Y(
        OR4_260_Y));
    OR4 OR4_567 (.A(\R_DATA_TEMPR8[39] ), .B(\R_DATA_TEMPR9[39] ), .C(
        \R_DATA_TEMPR10[39] ), .D(\R_DATA_TEMPR11[39] ), .Y(OR4_567_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%9%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R9C0 (.A_DOUT({
        \R_DATA_TEMPR9[39] , \R_DATA_TEMPR9[38] , \R_DATA_TEMPR9[37] , 
        \R_DATA_TEMPR9[36] , \R_DATA_TEMPR9[35] , \R_DATA_TEMPR9[34] , 
        \R_DATA_TEMPR9[33] , \R_DATA_TEMPR9[32] , \R_DATA_TEMPR9[31] , 
        \R_DATA_TEMPR9[30] , \R_DATA_TEMPR9[29] , \R_DATA_TEMPR9[28] , 
        \R_DATA_TEMPR9[27] , \R_DATA_TEMPR9[26] , \R_DATA_TEMPR9[25] , 
        \R_DATA_TEMPR9[24] , \R_DATA_TEMPR9[23] , \R_DATA_TEMPR9[22] , 
        \R_DATA_TEMPR9[21] , \R_DATA_TEMPR9[20] }), .B_DOUT({
        \R_DATA_TEMPR9[19] , \R_DATA_TEMPR9[18] , \R_DATA_TEMPR9[17] , 
        \R_DATA_TEMPR9[16] , \R_DATA_TEMPR9[15] , \R_DATA_TEMPR9[14] , 
        \R_DATA_TEMPR9[13] , \R_DATA_TEMPR9[12] , \R_DATA_TEMPR9[11] , 
        \R_DATA_TEMPR9[10] , \R_DATA_TEMPR9[9] , \R_DATA_TEMPR9[8] , 
        \R_DATA_TEMPR9[7] , \R_DATA_TEMPR9[6] , \R_DATA_TEMPR9[5] , 
        \R_DATA_TEMPR9[4] , \R_DATA_TEMPR9[3] , \R_DATA_TEMPR9[2] , 
        \R_DATA_TEMPR9[1] , \R_DATA_TEMPR9[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[9][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[2] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_406 (.A(\R_DATA_TEMPR36[17] ), .B(\R_DATA_TEMPR37[17] ), 
        .C(\R_DATA_TEMPR38[17] ), .D(\R_DATA_TEMPR39[17] ), .Y(
        OR4_406_Y));
    OR4 OR4_443 (.A(\R_DATA_TEMPR12[38] ), .B(\R_DATA_TEMPR13[38] ), 
        .C(\R_DATA_TEMPR14[38] ), .D(\R_DATA_TEMPR15[38] ), .Y(
        OR4_443_Y));
    OR4 OR4_669 (.A(\R_DATA_TEMPR24[20] ), .B(\R_DATA_TEMPR25[20] ), 
        .C(\R_DATA_TEMPR26[20] ), .D(\R_DATA_TEMPR27[20] ), .Y(
        OR4_669_Y));
    OR4 OR4_641 (.A(\R_DATA_TEMPR44[16] ), .B(\R_DATA_TEMPR45[16] ), 
        .C(\R_DATA_TEMPR46[16] ), .D(\R_DATA_TEMPR47[16] ), .Y(
        OR4_641_Y));
    OR4 OR4_184 (.A(\R_DATA_TEMPR20[15] ), .B(\R_DATA_TEMPR21[15] ), 
        .C(\R_DATA_TEMPR22[15] ), .D(\R_DATA_TEMPR23[15] ), .Y(
        OR4_184_Y));
    OR4 OR4_311 (.A(\R_DATA_TEMPR36[38] ), .B(\R_DATA_TEMPR37[38] ), 
        .C(\R_DATA_TEMPR38[38] ), .D(\R_DATA_TEMPR39[38] ), .Y(
        OR4_311_Y));
    OR4 OR4_476 (.A(\R_DATA_TEMPR28[24] ), .B(\R_DATA_TEMPR29[24] ), 
        .C(\R_DATA_TEMPR30[24] ), .D(\R_DATA_TEMPR31[24] ), .Y(
        OR4_476_Y));
    OR4 OR4_248 (.A(\R_DATA_TEMPR36[35] ), .B(\R_DATA_TEMPR37[35] ), 
        .C(\R_DATA_TEMPR38[35] ), .D(\R_DATA_TEMPR39[35] ), .Y(
        OR4_248_Y));
    OR4 OR4_757 (.A(OR4_635_Y), .B(OR4_798_Y), .C(OR4_82_Y), .D(
        OR4_674_Y), .Y(OR4_757_Y));
    OR4 OR4_754 (.A(\R_DATA_TEMPR56[15] ), .B(\R_DATA_TEMPR57[15] ), 
        .C(\R_DATA_TEMPR58[15] ), .D(\R_DATA_TEMPR59[15] ), .Y(
        OR4_754_Y));
    OR4 OR4_302 (.A(\R_DATA_TEMPR60[16] ), .B(\R_DATA_TEMPR61[16] ), 
        .C(\R_DATA_TEMPR62[16] ), .D(\R_DATA_TEMPR63[16] ), .Y(
        OR4_302_Y));
    OR4 OR4_266 (.A(OR4_418_Y), .B(OR4_119_Y), .C(OR4_385_Y), .D(
        OR4_613_Y), .Y(OR4_266_Y));
    OR4 OR4_10 (.A(\R_DATA_TEMPR56[37] ), .B(\R_DATA_TEMPR57[37] ), .C(
        \R_DATA_TEMPR58[37] ), .D(\R_DATA_TEMPR59[37] ), .Y(OR4_10_Y));
    OR4 OR4_25 (.A(\R_DATA_TEMPR60[25] ), .B(\R_DATA_TEMPR61[25] ), .C(
        \R_DATA_TEMPR62[25] ), .D(\R_DATA_TEMPR63[25] ), .Y(OR4_25_Y));
    OR4 OR4_76 (.A(\R_DATA_TEMPR56[28] ), .B(\R_DATA_TEMPR57[28] ), .C(
        \R_DATA_TEMPR58[28] ), .D(\R_DATA_TEMPR59[28] ), .Y(OR4_76_Y));
    OR4 OR4_410 (.A(\R_DATA_TEMPR4[11] ), .B(\R_DATA_TEMPR5[11] ), .C(
        \R_DATA_TEMPR6[11] ), .D(\R_DATA_TEMPR7[11] ), .Y(OR4_410_Y));
    OR4 OR4_339 (.A(\R_DATA_TEMPR24[34] ), .B(\R_DATA_TEMPR25[34] ), 
        .C(\R_DATA_TEMPR26[34] ), .D(\R_DATA_TEMPR27[34] ), .Y(
        OR4_339_Y));
    OR4 OR4_193 (.A(OR4_378_Y), .B(OR4_766_Y), .C(OR4_747_Y), .D(
        OR4_597_Y), .Y(OR4_193_Y));
    OR4 OR4_372 (.A(\R_DATA_TEMPR56[29] ), .B(\R_DATA_TEMPR57[29] ), 
        .C(\R_DATA_TEMPR58[29] ), .D(\R_DATA_TEMPR59[29] ), .Y(
        OR4_372_Y));
    OR4 OR4_525 (.A(\R_DATA_TEMPR40[7] ), .B(\R_DATA_TEMPR41[7] ), .C(
        \R_DATA_TEMPR42[7] ), .D(\R_DATA_TEMPR43[7] ), .Y(OR4_525_Y));
    OR4 OR4_17 (.A(\R_DATA_TEMPR12[1] ), .B(\R_DATA_TEMPR13[1] ), .C(
        \R_DATA_TEMPR14[1] ), .D(\R_DATA_TEMPR15[1] ), .Y(OR4_17_Y));
    OR4 OR4_781 (.A(\R_DATA_TEMPR12[0] ), .B(\R_DATA_TEMPR13[0] ), .C(
        \R_DATA_TEMPR14[0] ), .D(\R_DATA_TEMPR15[0] ), .Y(OR4_781_Y));
    OR4 OR4_664 (.A(OR4_199_Y), .B(OR4_323_Y), .C(OR4_414_Y), .D(
        OR4_789_Y), .Y(OR4_664_Y));
    CFG3 #( .INIT(8'h20) )  CFG3_14 (.A(W_ADDR[13]), .B(W_ADDR[12]), 
        .C(W_ADDR[11]), .Y(CFG3_14_Y));
    OR4 OR4_623 (.A(OR4_645_Y), .B(OR4_515_Y), .C(OR4_372_Y), .D(
        OR4_626_Y), .Y(OR4_623_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%4%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R4C0 (.A_DOUT({
        \R_DATA_TEMPR4[39] , \R_DATA_TEMPR4[38] , \R_DATA_TEMPR4[37] , 
        \R_DATA_TEMPR4[36] , \R_DATA_TEMPR4[35] , \R_DATA_TEMPR4[34] , 
        \R_DATA_TEMPR4[33] , \R_DATA_TEMPR4[32] , \R_DATA_TEMPR4[31] , 
        \R_DATA_TEMPR4[30] , \R_DATA_TEMPR4[29] , \R_DATA_TEMPR4[28] , 
        \R_DATA_TEMPR4[27] , \R_DATA_TEMPR4[26] , \R_DATA_TEMPR4[25] , 
        \R_DATA_TEMPR4[24] , \R_DATA_TEMPR4[23] , \R_DATA_TEMPR4[22] , 
        \R_DATA_TEMPR4[21] , \R_DATA_TEMPR4[20] }), .B_DOUT({
        \R_DATA_TEMPR4[19] , \R_DATA_TEMPR4[18] , \R_DATA_TEMPR4[17] , 
        \R_DATA_TEMPR4[16] , \R_DATA_TEMPR4[15] , \R_DATA_TEMPR4[14] , 
        \R_DATA_TEMPR4[13] , \R_DATA_TEMPR4[12] , \R_DATA_TEMPR4[11] , 
        \R_DATA_TEMPR4[10] , \R_DATA_TEMPR4[9] , \R_DATA_TEMPR4[8] , 
        \R_DATA_TEMPR4[7] , \R_DATA_TEMPR4[6] , \R_DATA_TEMPR4[5] , 
        \R_DATA_TEMPR4[4] , \R_DATA_TEMPR4[3] , \R_DATA_TEMPR4[2] , 
        \R_DATA_TEMPR4[1] , \R_DATA_TEMPR4[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[4][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[1] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_586 (.A(OR4_790_Y), .B(OR4_127_Y), .C(OR4_262_Y), .D(
        OR4_156_Y), .Y(OR4_586_Y));
    OR4 OR4_200 (.A(\R_DATA_TEMPR36[14] ), .B(\R_DATA_TEMPR37[14] ), 
        .C(\R_DATA_TEMPR38[14] ), .D(\R_DATA_TEMPR39[14] ), .Y(
        OR4_200_Y));
    OR4 OR4_507 (.A(OR4_308_Y), .B(OR4_452_Y), .C(OR4_183_Y), .D(
        OR4_604_Y), .Y(OR4_507_Y));
    OR4 OR4_270 (.A(OR4_792_Y), .B(OR4_130_Y), .C(OR4_671_Y), .D(
        OR4_296_Y), .Y(OR4_270_Y));
    OR4 OR4_577 (.A(\R_DATA_TEMPR52[38] ), .B(\R_DATA_TEMPR53[38] ), 
        .C(\R_DATA_TEMPR54[38] ), .D(\R_DATA_TEMPR55[38] ), .Y(
        OR4_577_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[12]  (.A(CFG3_11_Y), .B(
        CFG2_1_Y), .Y(\BLKY2[12] ));
    OR4 OR4_739 (.A(\R_DATA_TEMPR40[35] ), .B(\R_DATA_TEMPR41[35] ), 
        .C(\R_DATA_TEMPR42[35] ), .D(\R_DATA_TEMPR43[35] ), .Y(
        OR4_739_Y));
    OR4 OR4_541 (.A(\R_DATA_TEMPR12[11] ), .B(\R_DATA_TEMPR13[11] ), 
        .C(\R_DATA_TEMPR14[11] ), .D(\R_DATA_TEMPR15[11] ), .Y(
        OR4_541_Y));
    OR4 OR4_192 (.A(\R_DATA_TEMPR12[6] ), .B(\R_DATA_TEMPR13[6] ), .C(
        \R_DATA_TEMPR14[6] ), .D(\R_DATA_TEMPR15[6] ), .Y(OR4_192_Y));
    OR4 OR4_319 (.A(\R_DATA_TEMPR40[18] ), .B(\R_DATA_TEMPR41[18] ), 
        .C(\R_DATA_TEMPR42[18] ), .D(\R_DATA_TEMPR43[18] ), .Y(
        OR4_319_Y));
    OR4 OR4_609 (.A(\R_DATA_TEMPR36[23] ), .B(\R_DATA_TEMPR37[23] ), 
        .C(\R_DATA_TEMPR38[23] ), .D(\R_DATA_TEMPR39[23] ), .Y(
        OR4_609_Y));
    OR4 OR4_123 (.A(OR4_365_Y), .B(OR4_640_Y), .C(OR4_566_Y), .D(
        OR4_247_Y), .Y(OR4_123_Y));
    OR4 OR4_679 (.A(\R_DATA_TEMPR48[4] ), .B(\R_DATA_TEMPR49[4] ), .C(
        \R_DATA_TEMPR50[4] ), .D(\R_DATA_TEMPR51[4] ), .Y(OR4_679_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[2]  (.A(CFG3_8_Y), .B(CFG2_2_Y), 
        .Y(\BLKX2[2] ));
    OR4 OR4_206 (.A(\R_DATA_TEMPR28[23] ), .B(\R_DATA_TEMPR29[23] ), 
        .C(\R_DATA_TEMPR30[23] ), .D(\R_DATA_TEMPR31[23] ), .Y(
        OR4_206_Y));
    OR4 OR4_533 (.A(OR4_20_Y), .B(OR4_177_Y), .C(OR4_704_Y), .D(
        OR4_324_Y), .Y(OR4_533_Y));
    CFG2 #( .INIT(4'h8) )  CFG2_1 (.A(R_EN), .B(R_ADDR[14]), .Y(
        CFG2_1_Y));
    OR4 OR4_70 (.A(\R_DATA_TEMPR28[30] ), .B(\R_DATA_TEMPR29[30] ), .C(
        \R_DATA_TEMPR30[30] ), .D(\R_DATA_TEMPR31[30] ), .Y(OR4_70_Y));
    OR4 OR4_588 (.A(\R_DATA_TEMPR24[22] ), .B(\R_DATA_TEMPR25[22] ), 
        .C(\R_DATA_TEMPR26[22] ), .D(\R_DATA_TEMPR27[22] ), .Y(
        OR4_588_Y));
    OR4 OR4_58 (.A(\R_DATA_TEMPR20[12] ), .B(\R_DATA_TEMPR21[12] ), .C(
        \R_DATA_TEMPR22[12] ), .D(\R_DATA_TEMPR23[12] ), .Y(OR4_58_Y));
    OR4 OR4_276 (.A(\R_DATA_TEMPR44[34] ), .B(\R_DATA_TEMPR45[34] ), 
        .C(\R_DATA_TEMPR46[34] ), .D(\R_DATA_TEMPR47[34] ), .Y(
        OR4_276_Y));
    OR4 OR4_242 (.A(\R_DATA_TEMPR24[14] ), .B(\R_DATA_TEMPR25[14] ), 
        .C(\R_DATA_TEMPR26[14] ), .D(\R_DATA_TEMPR27[14] ), .Y(
        OR4_242_Y));
    OR4 OR4_77 (.A(OR4_211_Y), .B(OR4_488_Y), .C(OR4_67_Y), .D(
        OR4_205_Y), .Y(OR4_77_Y));
    OR4 OR4_604 (.A(\R_DATA_TEMPR44[5] ), .B(\R_DATA_TEMPR45[5] ), .C(
        \R_DATA_TEMPR46[5] ), .D(\R_DATA_TEMPR47[5] ), .Y(OR4_604_Y));
    OR4 OR4_299 (.A(\R_DATA_TEMPR20[11] ), .B(\R_DATA_TEMPR21[11] ), 
        .C(\R_DATA_TEMPR22[11] ), .D(\R_DATA_TEMPR23[11] ), .Y(
        OR4_299_Y));
    OR4 OR4_674 (.A(\R_DATA_TEMPR12[14] ), .B(\R_DATA_TEMPR13[14] ), 
        .C(\R_DATA_TEMPR14[14] ), .D(\R_DATA_TEMPR15[14] ), .Y(
        OR4_674_Y));
    OR4 OR4_455 (.A(\R_DATA_TEMPR40[8] ), .B(\R_DATA_TEMPR41[8] ), .C(
        \R_DATA_TEMPR42[8] ), .D(\R_DATA_TEMPR43[8] ), .Y(OR4_455_Y));
    OR4 OR4_486 (.A(\R_DATA_TEMPR52[13] ), .B(\R_DATA_TEMPR53[13] ), 
        .C(\R_DATA_TEMPR54[13] ), .D(\R_DATA_TEMPR55[13] ), .Y(
        OR4_486_Y));
    OR4 \OR4_R_DATA[5]  (.A(OR4_123_Y), .B(OR4_759_Y), .C(OR4_507_Y), 
        .D(OR4_664_Y), .Y(R_DATA[5]));
    OR4 OR4_340 (.A(\R_DATA_TEMPR8[21] ), .B(\R_DATA_TEMPR9[21] ), .C(
        \R_DATA_TEMPR10[21] ), .D(\R_DATA_TEMPR11[21] ), .Y(OR4_340_Y));
    OR4 OR4_719 (.A(\R_DATA_TEMPR56[10] ), .B(\R_DATA_TEMPR57[10] ), 
        .C(\R_DATA_TEMPR58[10] ), .D(\R_DATA_TEMPR59[10] ), .Y(
        OR4_719_Y));
    OR4 \OR4_R_DATA[11]  (.A(OR4_0_Y), .B(OR4_765_Y), .C(OR4_785_Y), 
        .D(OR4_534_Y), .Y(R_DATA[11]));
    OR4 OR4_122 (.A(\R_DATA_TEMPR24[1] ), .B(\R_DATA_TEMPR25[1] ), .C(
        \R_DATA_TEMPR26[1] ), .D(\R_DATA_TEMPR27[1] ), .Y(OR4_122_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R44C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%44%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R44C0 (
        .A_DOUT({\R_DATA_TEMPR44[39] , \R_DATA_TEMPR44[38] , 
        \R_DATA_TEMPR44[37] , \R_DATA_TEMPR44[36] , 
        \R_DATA_TEMPR44[35] , \R_DATA_TEMPR44[34] , 
        \R_DATA_TEMPR44[33] , \R_DATA_TEMPR44[32] , 
        \R_DATA_TEMPR44[31] , \R_DATA_TEMPR44[30] , 
        \R_DATA_TEMPR44[29] , \R_DATA_TEMPR44[28] , 
        \R_DATA_TEMPR44[27] , \R_DATA_TEMPR44[26] , 
        \R_DATA_TEMPR44[25] , \R_DATA_TEMPR44[24] , 
        \R_DATA_TEMPR44[23] , \R_DATA_TEMPR44[22] , 
        \R_DATA_TEMPR44[21] , \R_DATA_TEMPR44[20] }), .B_DOUT({
        \R_DATA_TEMPR44[19] , \R_DATA_TEMPR44[18] , 
        \R_DATA_TEMPR44[17] , \R_DATA_TEMPR44[16] , 
        \R_DATA_TEMPR44[15] , \R_DATA_TEMPR44[14] , 
        \R_DATA_TEMPR44[13] , \R_DATA_TEMPR44[12] , 
        \R_DATA_TEMPR44[11] , \R_DATA_TEMPR44[10] , 
        \R_DATA_TEMPR44[9] , \R_DATA_TEMPR44[8] , \R_DATA_TEMPR44[7] , 
        \R_DATA_TEMPR44[6] , \R_DATA_TEMPR44[5] , \R_DATA_TEMPR44[4] , 
        \R_DATA_TEMPR44[3] , \R_DATA_TEMPR44[2] , \R_DATA_TEMPR44[1] , 
        \R_DATA_TEMPR44[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[44][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[11] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[11] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_382 (.A(\R_DATA_TEMPR52[3] ), .B(\R_DATA_TEMPR53[3] ), .C(
        \R_DATA_TEMPR54[3] ), .D(\R_DATA_TEMPR55[3] ), .Y(OR4_382_Y));
    OR4 \OR4_R_DATA[9]  (.A(OR4_101_Y), .B(OR4_266_Y), .C(OR4_460_Y), 
        .D(OR4_620_Y), .Y(R_DATA[9]));
    OR4 OR4_18 (.A(OR4_166_Y), .B(OR4_35_Y), .C(OR4_699_Y), .D(
        OR4_306_Y), .Y(OR4_18_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R35C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%35%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R35C0 (
        .A_DOUT({\R_DATA_TEMPR35[39] , \R_DATA_TEMPR35[38] , 
        \R_DATA_TEMPR35[37] , \R_DATA_TEMPR35[36] , 
        \R_DATA_TEMPR35[35] , \R_DATA_TEMPR35[34] , 
        \R_DATA_TEMPR35[33] , \R_DATA_TEMPR35[32] , 
        \R_DATA_TEMPR35[31] , \R_DATA_TEMPR35[30] , 
        \R_DATA_TEMPR35[29] , \R_DATA_TEMPR35[28] , 
        \R_DATA_TEMPR35[27] , \R_DATA_TEMPR35[26] , 
        \R_DATA_TEMPR35[25] , \R_DATA_TEMPR35[24] , 
        \R_DATA_TEMPR35[23] , \R_DATA_TEMPR35[22] , 
        \R_DATA_TEMPR35[21] , \R_DATA_TEMPR35[20] }), .B_DOUT({
        \R_DATA_TEMPR35[19] , \R_DATA_TEMPR35[18] , 
        \R_DATA_TEMPR35[17] , \R_DATA_TEMPR35[16] , 
        \R_DATA_TEMPR35[15] , \R_DATA_TEMPR35[14] , 
        \R_DATA_TEMPR35[13] , \R_DATA_TEMPR35[12] , 
        \R_DATA_TEMPR35[11] , \R_DATA_TEMPR35[10] , 
        \R_DATA_TEMPR35[9] , \R_DATA_TEMPR35[8] , \R_DATA_TEMPR35[7] , 
        \R_DATA_TEMPR35[6] , \R_DATA_TEMPR35[5] , \R_DATA_TEMPR35[4] , 
        \R_DATA_TEMPR35[3] , \R_DATA_TEMPR35[2] , \R_DATA_TEMPR35[1] , 
        \R_DATA_TEMPR35[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[35][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[8] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[8] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_513 (.A(\R_DATA_TEMPR12[4] ), .B(\R_DATA_TEMPR13[4] ), .C(
        \R_DATA_TEMPR14[4] ), .D(\R_DATA_TEMPR15[4] ), .Y(OR4_513_Y));
    OR4 OR4_34 (.A(\R_DATA_TEMPR32[0] ), .B(\R_DATA_TEMPR33[0] ), .C(
        \R_DATA_TEMPR34[0] ), .D(\R_DATA_TEMPR35[0] ), .Y(OR4_34_Y));
    OR4 OR4_454 (.A(\R_DATA_TEMPR48[16] ), .B(\R_DATA_TEMPR49[16] ), 
        .C(\R_DATA_TEMPR50[16] ), .D(\R_DATA_TEMPR51[16] ), .Y(
        OR4_454_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[11]  (.A(CFG3_12_Y), .B(
        CFG2_1_Y), .Y(\BLKY2[11] ));
    OR4 \OR4_R_DATA[35]  (.A(OR4_74_Y), .B(OR4_461_Y), .C(OR4_778_Y), 
        .D(OR4_545_Y), .Y(R_DATA[35]));
    OR4 \OR4_R_DATA[10]  (.A(OR4_655_Y), .B(OR4_33_Y), .C(OR4_398_Y), 
        .D(OR4_88_Y), .Y(R_DATA[10]));
    OR4 OR4_229 (.A(OR4_598_Y), .B(OR4_72_Y), .C(OR4_464_Y), .D(
        OR4_591_Y), .Y(OR4_229_Y));
    OR4 OR4_356 (.A(OR4_347_Y), .B(OR4_226_Y), .C(OR4_75_Y), .D(
        OR4_234_Y), .Y(OR4_356_Y));
    OR4 OR4_797 (.A(\R_DATA_TEMPR20[29] ), .B(\R_DATA_TEMPR21[29] ), 
        .C(\R_DATA_TEMPR22[29] ), .D(\R_DATA_TEMPR23[29] ), .Y(
        OR4_797_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R41C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%41%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R41C0 (
        .A_DOUT({\R_DATA_TEMPR41[39] , \R_DATA_TEMPR41[38] , 
        \R_DATA_TEMPR41[37] , \R_DATA_TEMPR41[36] , 
        \R_DATA_TEMPR41[35] , \R_DATA_TEMPR41[34] , 
        \R_DATA_TEMPR41[33] , \R_DATA_TEMPR41[32] , 
        \R_DATA_TEMPR41[31] , \R_DATA_TEMPR41[30] , 
        \R_DATA_TEMPR41[29] , \R_DATA_TEMPR41[28] , 
        \R_DATA_TEMPR41[27] , \R_DATA_TEMPR41[26] , 
        \R_DATA_TEMPR41[25] , \R_DATA_TEMPR41[24] , 
        \R_DATA_TEMPR41[23] , \R_DATA_TEMPR41[22] , 
        \R_DATA_TEMPR41[21] , \R_DATA_TEMPR41[20] }), .B_DOUT({
        \R_DATA_TEMPR41[19] , \R_DATA_TEMPR41[18] , 
        \R_DATA_TEMPR41[17] , \R_DATA_TEMPR41[16] , 
        \R_DATA_TEMPR41[15] , \R_DATA_TEMPR41[14] , 
        \R_DATA_TEMPR41[13] , \R_DATA_TEMPR41[12] , 
        \R_DATA_TEMPR41[11] , \R_DATA_TEMPR41[10] , 
        \R_DATA_TEMPR41[9] , \R_DATA_TEMPR41[8] , \R_DATA_TEMPR41[7] , 
        \R_DATA_TEMPR41[6] , \R_DATA_TEMPR41[5] , \R_DATA_TEMPR41[4] , 
        \R_DATA_TEMPR41[3] , \R_DATA_TEMPR41[2] , \R_DATA_TEMPR41[1] , 
        \R_DATA_TEMPR41[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[41][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[10] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[10] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_794 (.A(\R_DATA_TEMPR36[7] ), .B(\R_DATA_TEMPR37[7] ), .C(
        \R_DATA_TEMPR38[7] ), .D(\R_DATA_TEMPR39[7] ), .Y(OR4_794_Y));
    OR4 OR4_261 (.A(\R_DATA_TEMPR48[6] ), .B(\R_DATA_TEMPR49[6] ), .C(
        \R_DATA_TEMPR50[6] ), .D(\R_DATA_TEMPR51[6] ), .Y(OR4_261_Y));
    OR4 OR4_29 (.A(\R_DATA_TEMPR28[17] ), .B(\R_DATA_TEMPR29[17] ), .C(
        \R_DATA_TEMPR30[17] ), .D(\R_DATA_TEMPR31[17] ), .Y(OR4_29_Y));
    OR4 \OR4_R_DATA[16]  (.A(OR4_373_Y), .B(OR4_6_Y), .C(OR4_149_Y), 
        .D(OR4_191_Y), .Y(R_DATA[16]));
    OR4 OR4_280 (.A(\R_DATA_TEMPR8[34] ), .B(\R_DATA_TEMPR9[34] ), .C(
        \R_DATA_TEMPR10[34] ), .D(\R_DATA_TEMPR11[34] ), .Y(OR4_280_Y));
    OR4 OR4_587 (.A(OR4_165_Y), .B(OR4_505_Y), .C(OR4_779_Y), .D(
        OR4_477_Y), .Y(OR4_587_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%23%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R23C0 (
        .A_DOUT({\R_DATA_TEMPR23[39] , \R_DATA_TEMPR23[38] , 
        \R_DATA_TEMPR23[37] , \R_DATA_TEMPR23[36] , 
        \R_DATA_TEMPR23[35] , \R_DATA_TEMPR23[34] , 
        \R_DATA_TEMPR23[33] , \R_DATA_TEMPR23[32] , 
        \R_DATA_TEMPR23[31] , \R_DATA_TEMPR23[30] , 
        \R_DATA_TEMPR23[29] , \R_DATA_TEMPR23[28] , 
        \R_DATA_TEMPR23[27] , \R_DATA_TEMPR23[26] , 
        \R_DATA_TEMPR23[25] , \R_DATA_TEMPR23[24] , 
        \R_DATA_TEMPR23[23] , \R_DATA_TEMPR23[22] , 
        \R_DATA_TEMPR23[21] , \R_DATA_TEMPR23[20] }), .B_DOUT({
        \R_DATA_TEMPR23[19] , \R_DATA_TEMPR23[18] , 
        \R_DATA_TEMPR23[17] , \R_DATA_TEMPR23[16] , 
        \R_DATA_TEMPR23[15] , \R_DATA_TEMPR23[14] , 
        \R_DATA_TEMPR23[13] , \R_DATA_TEMPR23[12] , 
        \R_DATA_TEMPR23[11] , \R_DATA_TEMPR23[10] , 
        \R_DATA_TEMPR23[9] , \R_DATA_TEMPR23[8] , \R_DATA_TEMPR23[7] , 
        \R_DATA_TEMPR23[6] , \R_DATA_TEMPR23[5] , \R_DATA_TEMPR23[4] , 
        \R_DATA_TEMPR23[3] , \R_DATA_TEMPR23[2] , \R_DATA_TEMPR23[1] , 
        \R_DATA_TEMPR23[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[5] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[5] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_545 (.A(OR4_753_Y), .B(OR4_519_Y), .C(OR4_543_Y), .D(
        OR4_672_Y), .Y(OR4_545_Y));
    OR4 OR4_233 (.A(\R_DATA_TEMPR28[31] ), .B(\R_DATA_TEMPR29[31] ), 
        .C(\R_DATA_TEMPR30[31] ), .D(\R_DATA_TEMPR31[31] ), .Y(
        OR4_233_Y));
    OR4 OR4_562 (.A(\R_DATA_TEMPR12[17] ), .B(\R_DATA_TEMPR13[17] ), 
        .C(\R_DATA_TEMPR14[17] ), .D(\R_DATA_TEMPR15[17] ), .Y(
        OR4_562_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%17%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R17C0 (
        .A_DOUT({\R_DATA_TEMPR17[39] , \R_DATA_TEMPR17[38] , 
        \R_DATA_TEMPR17[37] , \R_DATA_TEMPR17[36] , 
        \R_DATA_TEMPR17[35] , \R_DATA_TEMPR17[34] , 
        \R_DATA_TEMPR17[33] , \R_DATA_TEMPR17[32] , 
        \R_DATA_TEMPR17[31] , \R_DATA_TEMPR17[30] , 
        \R_DATA_TEMPR17[29] , \R_DATA_TEMPR17[28] , 
        \R_DATA_TEMPR17[27] , \R_DATA_TEMPR17[26] , 
        \R_DATA_TEMPR17[25] , \R_DATA_TEMPR17[24] , 
        \R_DATA_TEMPR17[23] , \R_DATA_TEMPR17[22] , 
        \R_DATA_TEMPR17[21] , \R_DATA_TEMPR17[20] }), .B_DOUT({
        \R_DATA_TEMPR17[19] , \R_DATA_TEMPR17[18] , 
        \R_DATA_TEMPR17[17] , \R_DATA_TEMPR17[16] , 
        \R_DATA_TEMPR17[15] , \R_DATA_TEMPR17[14] , 
        \R_DATA_TEMPR17[13] , \R_DATA_TEMPR17[12] , 
        \R_DATA_TEMPR17[11] , \R_DATA_TEMPR17[10] , 
        \R_DATA_TEMPR17[9] , \R_DATA_TEMPR17[8] , \R_DATA_TEMPR17[7] , 
        \R_DATA_TEMPR17[6] , \R_DATA_TEMPR17[5] , \R_DATA_TEMPR17[4] , 
        \R_DATA_TEMPR17[3] , \R_DATA_TEMPR17[2] , \R_DATA_TEMPR17[1] , 
        \R_DATA_TEMPR17[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[4] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_689 (.A(OR4_2_Y), .B(OR4_295_Y), .C(OR4_676_Y), .D(
        OR4_796_Y), .Y(OR4_689_Y));
    OR4 OR4_643 (.A(\R_DATA_TEMPR12[26] ), .B(\R_DATA_TEMPR13[26] ), 
        .C(\R_DATA_TEMPR14[26] ), .D(\R_DATA_TEMPR15[26] ), .Y(
        OR4_643_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[4]  (.A(CFG3_11_Y), .B(CFG2_0_Y)
        , .Y(\BLKY2[4] ));
    OR4 OR4_286 (.A(\R_DATA_TEMPR24[11] ), .B(\R_DATA_TEMPR25[11] ), 
        .C(\R_DATA_TEMPR26[11] ), .D(\R_DATA_TEMPR27[11] ), .Y(
        OR4_286_Y));
    OR4 OR4_78 (.A(\R_DATA_TEMPR44[29] ), .B(\R_DATA_TEMPR45[29] ), .C(
        \R_DATA_TEMPR46[29] ), .D(\R_DATA_TEMPR47[29] ), .Y(OR4_78_Y));
    OR4 \OR4_R_DATA[8]  (.A(OR4_402_Y), .B(OR4_492_Y), .C(OR4_303_Y), 
        .D(OR4_599_Y), .Y(R_DATA[8]));
    OR4 OR4_564 (.A(\R_DATA_TEMPR60[13] ), .B(\R_DATA_TEMPR61[13] ), 
        .C(\R_DATA_TEMPR62[13] ), .D(\R_DATA_TEMPR63[13] ), .Y(
        OR4_564_Y));
    OR4 OR4_154 (.A(\R_DATA_TEMPR52[25] ), .B(\R_DATA_TEMPR53[25] ), 
        .C(\R_DATA_TEMPR54[25] ), .D(\R_DATA_TEMPR55[25] ), .Y(
        OR4_154_Y));
    OR4 OR4_727 (.A(\R_DATA_TEMPR40[16] ), .B(\R_DATA_TEMPR41[16] ), 
        .C(\R_DATA_TEMPR42[16] ), .D(\R_DATA_TEMPR43[16] ), .Y(
        OR4_727_Y));
    OR4 OR4_684 (.A(\R_DATA_TEMPR56[8] ), .B(\R_DATA_TEMPR57[8] ), .C(
        \R_DATA_TEMPR58[8] ), .D(\R_DATA_TEMPR59[8] ), .Y(OR4_684_Y));
    OR4 OR4_724 (.A(\R_DATA_TEMPR36[8] ), .B(\R_DATA_TEMPR37[8] ), .C(
        \R_DATA_TEMPR38[8] ), .D(\R_DATA_TEMPR39[8] ), .Y(OR4_724_Y));
    OR4 OR4_638 (.A(\R_DATA_TEMPR24[39] ), .B(\R_DATA_TEMPR25[39] ), 
        .C(\R_DATA_TEMPR26[39] ), .D(\R_DATA_TEMPR27[39] ), .Y(
        OR4_638_Y));
    OR4 OR4_22 (.A(OR4_337_Y), .B(OR4_489_Y), .C(OR4_614_Y), .D(
        OR4_518_Y), .Y(OR4_22_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[15]  (.A(CFG3_13_Y), .B(
        CFG2_1_Y), .Y(\BLKY2[15] ));
    OR4 OR4_143 (.A(\R_DATA_TEMPR60[18] ), .B(\R_DATA_TEMPR61[18] ), 
        .C(\R_DATA_TEMPR62[18] ), .D(\R_DATA_TEMPR63[18] ), .Y(
        OR4_143_Y));
    OR4 OR4_632 (.A(\R_DATA_TEMPR20[4] ), .B(\R_DATA_TEMPR21[4] ), .C(
        \R_DATA_TEMPR22[4] ), .D(\R_DATA_TEMPR23[4] ), .Y(OR4_632_Y));
    OR4 OR4_213 (.A(\R_DATA_TEMPR32[32] ), .B(\R_DATA_TEMPR33[32] ), 
        .C(\R_DATA_TEMPR34[32] ), .D(\R_DATA_TEMPR35[32] ), .Y(
        OR4_213_Y));
    OR4 OR4_201 (.A(\R_DATA_TEMPR16[11] ), .B(\R_DATA_TEMPR17[11] ), 
        .C(\R_DATA_TEMPR18[11] ), .D(\R_DATA_TEMPR19[11] ), .Y(
        OR4_201_Y));
    OR4 OR4_361 (.A(\R_DATA_TEMPR16[29] ), .B(\R_DATA_TEMPR17[29] ), 
        .C(\R_DATA_TEMPR18[29] ), .D(\R_DATA_TEMPR19[29] ), .Y(
        OR4_361_Y));
    OR4 OR4_751 (.A(OR4_85_Y), .B(OR4_371_Y), .C(OR4_750_Y), .D(
        OR4_78_Y), .Y(OR4_751_Y));
    OR4 OR4_6 (.A(OR4_198_Y), .B(OR4_665_Y), .C(OR4_653_Y), .D(
        OR4_235_Y), .Y(OR4_6_Y));
    OR4 OR4_271 (.A(\R_DATA_TEMPR48[3] ), .B(\R_DATA_TEMPR49[3] ), .C(
        \R_DATA_TEMPR50[3] ), .D(\R_DATA_TEMPR51[3] ), .Y(OR4_271_Y));
    OR4 OR4_460 (.A(OR4_290_Y), .B(OR4_435_Y), .C(OR4_164_Y), .D(
        OR4_579_Y), .Y(OR4_460_Y));
    OR4 OR4_502 (.A(\R_DATA_TEMPR4[3] ), .B(\R_DATA_TEMPR5[3] ), .C(
        \R_DATA_TEMPR6[3] ), .D(\R_DATA_TEMPR7[3] ), .Y(OR4_502_Y));
    OR4 OR4_556 (.A(OR4_138_Y), .B(OR4_705_Y), .C(OR4_738_Y), .D(
        OR4_86_Y), .Y(OR4_556_Y));
    OR4 OR4_495 (.A(\R_DATA_TEMPR8[26] ), .B(\R_DATA_TEMPR9[26] ), .C(
        \R_DATA_TEMPR10[26] ), .D(\R_DATA_TEMPR11[26] ), .Y(OR4_495_Y));
    OR4 OR4_572 (.A(\R_DATA_TEMPR8[0] ), .B(\R_DATA_TEMPR9[0] ), .C(
        \R_DATA_TEMPR10[0] ), .D(\R_DATA_TEMPR11[0] ), .Y(OR4_572_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%3%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R3C0 (.A_DOUT({
        \R_DATA_TEMPR3[39] , \R_DATA_TEMPR3[38] , \R_DATA_TEMPR3[37] , 
        \R_DATA_TEMPR3[36] , \R_DATA_TEMPR3[35] , \R_DATA_TEMPR3[34] , 
        \R_DATA_TEMPR3[33] , \R_DATA_TEMPR3[32] , \R_DATA_TEMPR3[31] , 
        \R_DATA_TEMPR3[30] , \R_DATA_TEMPR3[29] , \R_DATA_TEMPR3[28] , 
        \R_DATA_TEMPR3[27] , \R_DATA_TEMPR3[26] , \R_DATA_TEMPR3[25] , 
        \R_DATA_TEMPR3[24] , \R_DATA_TEMPR3[23] , \R_DATA_TEMPR3[22] , 
        \R_DATA_TEMPR3[21] , \R_DATA_TEMPR3[20] }), .B_DOUT({
        \R_DATA_TEMPR3[19] , \R_DATA_TEMPR3[18] , \R_DATA_TEMPR3[17] , 
        \R_DATA_TEMPR3[16] , \R_DATA_TEMPR3[15] , \R_DATA_TEMPR3[14] , 
        \R_DATA_TEMPR3[13] , \R_DATA_TEMPR3[12] , \R_DATA_TEMPR3[11] , 
        \R_DATA_TEMPR3[10] , \R_DATA_TEMPR3[9] , \R_DATA_TEMPR3[8] , 
        \R_DATA_TEMPR3[7] , \R_DATA_TEMPR3[6] , \R_DATA_TEMPR3[5] , 
        \R_DATA_TEMPR3[4] , \R_DATA_TEMPR3[3] , \R_DATA_TEMPR3[2] , 
        \R_DATA_TEMPR3[1] , \R_DATA_TEMPR3[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[3][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_618 (.A(OR4_92_Y), .B(OR4_245_Y), .C(OR4_97_Y), .D(
        OR4_513_Y), .Y(OR4_618_Y));
    CFG3 #( .INIT(8'h4) )  CFG3_8 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_8_Y));
    OR4 \OR4_R_DATA[17]  (.A(OR4_170_Y), .B(OR4_552_Y), .C(OR4_752_Y), 
        .D(OR4_31_Y), .Y(R_DATA[17]));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[0]  (.A(CFG3_10_Y), .B(CFG2_0_Y)
        , .Y(\BLKY2[0] ));
    OR4 OR4_142 (.A(\R_DATA_TEMPR0[25] ), .B(\R_DATA_TEMPR1[25] ), .C(
        \R_DATA_TEMPR2[25] ), .D(\R_DATA_TEMPR3[25] ), .Y(OR4_142_Y));
    OR4 OR4_612 (.A(\R_DATA_TEMPR56[23] ), .B(\R_DATA_TEMPR57[23] ), 
        .C(\R_DATA_TEMPR58[23] ), .D(\R_DATA_TEMPR59[23] ), .Y(
        OR4_612_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R53C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%53%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R53C0 (
        .A_DOUT({\R_DATA_TEMPR53[39] , \R_DATA_TEMPR53[38] , 
        \R_DATA_TEMPR53[37] , \R_DATA_TEMPR53[36] , 
        \R_DATA_TEMPR53[35] , \R_DATA_TEMPR53[34] , 
        \R_DATA_TEMPR53[33] , \R_DATA_TEMPR53[32] , 
        \R_DATA_TEMPR53[31] , \R_DATA_TEMPR53[30] , 
        \R_DATA_TEMPR53[29] , \R_DATA_TEMPR53[28] , 
        \R_DATA_TEMPR53[27] , \R_DATA_TEMPR53[26] , 
        \R_DATA_TEMPR53[25] , \R_DATA_TEMPR53[24] , 
        \R_DATA_TEMPR53[23] , \R_DATA_TEMPR53[22] , 
        \R_DATA_TEMPR53[21] , \R_DATA_TEMPR53[20] }), .B_DOUT({
        \R_DATA_TEMPR53[19] , \R_DATA_TEMPR53[18] , 
        \R_DATA_TEMPR53[17] , \R_DATA_TEMPR53[16] , 
        \R_DATA_TEMPR53[15] , \R_DATA_TEMPR53[14] , 
        \R_DATA_TEMPR53[13] , \R_DATA_TEMPR53[12] , 
        \R_DATA_TEMPR53[11] , \R_DATA_TEMPR53[10] , 
        \R_DATA_TEMPR53[9] , \R_DATA_TEMPR53[8] , \R_DATA_TEMPR53[7] , 
        \R_DATA_TEMPR53[6] , \R_DATA_TEMPR53[5] , \R_DATA_TEMPR53[4] , 
        \R_DATA_TEMPR53[3] , \R_DATA_TEMPR53[2] , \R_DATA_TEMPR53[1] , 
        \R_DATA_TEMPR53[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[53][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[13] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[13] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_504 (.A(\R_DATA_TEMPR20[24] ), .B(\R_DATA_TEMPR21[24] ), 
        .C(\R_DATA_TEMPR22[24] ), .D(\R_DATA_TEMPR23[24] ), .Y(
        OR4_504_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%28%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R28C0 (
        .A_DOUT({\R_DATA_TEMPR28[39] , \R_DATA_TEMPR28[38] , 
        \R_DATA_TEMPR28[37] , \R_DATA_TEMPR28[36] , 
        \R_DATA_TEMPR28[35] , \R_DATA_TEMPR28[34] , 
        \R_DATA_TEMPR28[33] , \R_DATA_TEMPR28[32] , 
        \R_DATA_TEMPR28[31] , \R_DATA_TEMPR28[30] , 
        \R_DATA_TEMPR28[29] , \R_DATA_TEMPR28[28] , 
        \R_DATA_TEMPR28[27] , \R_DATA_TEMPR28[26] , 
        \R_DATA_TEMPR28[25] , \R_DATA_TEMPR28[24] , 
        \R_DATA_TEMPR28[23] , \R_DATA_TEMPR28[22] , 
        \R_DATA_TEMPR28[21] , \R_DATA_TEMPR28[20] }), .B_DOUT({
        \R_DATA_TEMPR28[19] , \R_DATA_TEMPR28[18] , 
        \R_DATA_TEMPR28[17] , \R_DATA_TEMPR28[16] , 
        \R_DATA_TEMPR28[15] , \R_DATA_TEMPR28[14] , 
        \R_DATA_TEMPR28[13] , \R_DATA_TEMPR28[12] , 
        \R_DATA_TEMPR28[11] , \R_DATA_TEMPR28[10] , 
        \R_DATA_TEMPR28[9] , \R_DATA_TEMPR28[8] , \R_DATA_TEMPR28[7] , 
        \R_DATA_TEMPR28[6] , \R_DATA_TEMPR28[5] , \R_DATA_TEMPR28[4] , 
        \R_DATA_TEMPR28[3] , \R_DATA_TEMPR28[2] , \R_DATA_TEMPR28[1] , 
        \R_DATA_TEMPR28[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[7] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_574 (.A(\R_DATA_TEMPR52[34] ), .B(\R_DATA_TEMPR53[34] ), 
        .C(\R_DATA_TEMPR54[34] ), .D(\R_DATA_TEMPR55[34] ), .Y(
        OR4_574_Y));
    OR4 OR4_494 (.A(\R_DATA_TEMPR8[22] ), .B(\R_DATA_TEMPR9[22] ), .C(
        \R_DATA_TEMPR10[22] ), .D(\R_DATA_TEMPR11[22] ), .Y(OR4_494_Y));
    OR4 OR4_558 (.A(\R_DATA_TEMPR44[39] ), .B(\R_DATA_TEMPR45[39] ), 
        .C(\R_DATA_TEMPR46[39] ), .D(\R_DATA_TEMPR47[39] ), .Y(
        OR4_558_Y));
    OR4 OR4_55 (.A(\R_DATA_TEMPR48[31] ), .B(\R_DATA_TEMPR49[31] ), .C(
        \R_DATA_TEMPR50[31] ), .D(\R_DATA_TEMPR51[31] ), .Y(OR4_55_Y));
    OR4 OR4_369 (.A(\R_DATA_TEMPR4[6] ), .B(\R_DATA_TEMPR5[6] ), .C(
        \R_DATA_TEMPR6[6] ), .D(\R_DATA_TEMPR7[6] ), .Y(OR4_369_Y));
    OR4 OR4_301 (.A(OR4_291_Y), .B(OR4_154_Y), .C(OR4_15_Y), .D(
        OR4_25_Y), .Y(OR4_301_Y));
    OR4 OR4_396 (.A(\R_DATA_TEMPR52[32] ), .B(\R_DATA_TEMPR53[32] ), 
        .C(\R_DATA_TEMPR54[32] ), .D(\R_DATA_TEMPR55[32] ), .Y(
        OR4_396_Y));
    OR4 OR4_249 (.A(\R_DATA_TEMPR40[6] ), .B(\R_DATA_TEMPR41[6] ), .C(
        \R_DATA_TEMPR42[6] ), .D(\R_DATA_TEMPR43[6] ), .Y(OR4_249_Y));
    OR4 OR4_371 (.A(\R_DATA_TEMPR36[29] ), .B(\R_DATA_TEMPR37[29] ), 
        .C(\R_DATA_TEMPR38[29] ), .D(\R_DATA_TEMPR39[29] ), .Y(
        OR4_371_Y));
    OR4 OR4_425 (.A(OR4_687_Y), .B(OR4_530_Y), .C(OR4_517_Y), .D(
        OR4_208_Y), .Y(OR4_425_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%0%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R0C0 (.A_DOUT({
        \R_DATA_TEMPR0[39] , \R_DATA_TEMPR0[38] , \R_DATA_TEMPR0[37] , 
        \R_DATA_TEMPR0[36] , \R_DATA_TEMPR0[35] , \R_DATA_TEMPR0[34] , 
        \R_DATA_TEMPR0[33] , \R_DATA_TEMPR0[32] , \R_DATA_TEMPR0[31] , 
        \R_DATA_TEMPR0[30] , \R_DATA_TEMPR0[29] , \R_DATA_TEMPR0[28] , 
        \R_DATA_TEMPR0[27] , \R_DATA_TEMPR0[26] , \R_DATA_TEMPR0[25] , 
        \R_DATA_TEMPR0[24] , \R_DATA_TEMPR0[23] , \R_DATA_TEMPR0[22] , 
        \R_DATA_TEMPR0[21] , \R_DATA_TEMPR0[20] }), .B_DOUT({
        \R_DATA_TEMPR0[19] , \R_DATA_TEMPR0[18] , \R_DATA_TEMPR0[17] , 
        \R_DATA_TEMPR0[16] , \R_DATA_TEMPR0[15] , \R_DATA_TEMPR0[14] , 
        \R_DATA_TEMPR0[13] , \R_DATA_TEMPR0[12] , \R_DATA_TEMPR0[11] , 
        \R_DATA_TEMPR0[10] , \R_DATA_TEMPR0[9] , \R_DATA_TEMPR0[8] , 
        \R_DATA_TEMPR0[7] , \R_DATA_TEMPR0[6] , \R_DATA_TEMPR0[5] , 
        \R_DATA_TEMPR0[4] , \R_DATA_TEMPR0[3] , \R_DATA_TEMPR0[2] , 
        \R_DATA_TEMPR0[1] , \R_DATA_TEMPR0[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[0][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_400 (.A(\R_DATA_TEMPR40[25] ), .B(\R_DATA_TEMPR41[25] ), 
        .C(\R_DATA_TEMPR42[25] ), .D(\R_DATA_TEMPR43[25] ), .Y(
        OR4_400_Y));
    OR4 OR4_636 (.A(\R_DATA_TEMPR0[0] ), .B(\R_DATA_TEMPR1[0] ), .C(
        \R_DATA_TEMPR2[0] ), .D(\R_DATA_TEMPR3[0] ), .Y(OR4_636_Y));
    OR4 \OR4_R_DATA[38]  (.A(OR4_144_Y), .B(OR4_37_Y), .C(OR4_472_Y), 
        .D(OR4_582_Y), .Y(R_DATA[38]));
    OR4 OR4_456 (.A(\R_DATA_TEMPR0[31] ), .B(\R_DATA_TEMPR1[31] ), .C(
        \R_DATA_TEMPR2[31] ), .D(\R_DATA_TEMPR3[31] ), .Y(OR4_456_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[5]  (.A(CFG3_6_Y), .B(CFG2_0_Y), 
        .Y(\BLKY2[5] ));
    OR4 OR4_470 (.A(\R_DATA_TEMPR24[3] ), .B(\R_DATA_TEMPR25[3] ), .C(
        \R_DATA_TEMPR26[3] ), .D(\R_DATA_TEMPR27[3] ), .Y(OR4_470_Y));
    OR4 OR4_352 (.A(\R_DATA_TEMPR4[18] ), .B(\R_DATA_TEMPR5[18] ), .C(
        \R_DATA_TEMPR6[18] ), .D(\R_DATA_TEMPR7[18] ), .Y(OR4_352_Y));
    OR4 OR4_15 (.A(\R_DATA_TEMPR56[25] ), .B(\R_DATA_TEMPR57[25] ), .C(
        \R_DATA_TEMPR58[25] ), .D(\R_DATA_TEMPR59[25] ), .Y(OR4_15_Y));
    OR4 OR4_424 (.A(\R_DATA_TEMPR4[10] ), .B(\R_DATA_TEMPR5[10] ), .C(
        \R_DATA_TEMPR6[10] ), .D(\R_DATA_TEMPR7[10] ), .Y(OR4_424_Y));
    OR4 OR4_281 (.A(\R_DATA_TEMPR12[13] ), .B(\R_DATA_TEMPR13[13] ), 
        .C(\R_DATA_TEMPR14[13] ), .D(\R_DATA_TEMPR15[13] ), .Y(
        OR4_281_Y));
    OR4 OR4_769 (.A(\R_DATA_TEMPR8[33] ), .B(\R_DATA_TEMPR9[33] ), .C(
        \R_DATA_TEMPR10[33] ), .D(\R_DATA_TEMPR11[33] ), .Y(OR4_769_Y));
    OR4 OR4_194 (.A(OR4_244_Y), .B(OR4_502_Y), .C(OR4_703_Y), .D(
        OR4_277_Y), .Y(OR4_194_Y));
    OR4 OR4_326 (.A(\R_DATA_TEMPR20[22] ), .B(\R_DATA_TEMPR21[22] ), 
        .C(\R_DATA_TEMPR22[22] ), .D(\R_DATA_TEMPR23[22] ), .Y(
        OR4_326_Y));
    OR4 OR4_747 (.A(\R_DATA_TEMPR24[36] ), .B(\R_DATA_TEMPR25[36] ), 
        .C(\R_DATA_TEMPR26[36] ), .D(\R_DATA_TEMPR27[36] ), .Y(
        OR4_747_Y));
    OR4 OR4_563 (.A(\R_DATA_TEMPR60[15] ), .B(\R_DATA_TEMPR61[15] ), 
        .C(\R_DATA_TEMPR62[15] ), .D(\R_DATA_TEMPR63[15] ), .Y(
        OR4_563_Y));
    OR4 OR4_93 (.A(\R_DATA_TEMPR12[22] ), .B(\R_DATA_TEMPR13[22] ), .C(
        \R_DATA_TEMPR14[22] ), .D(\R_DATA_TEMPR15[22] ), .Y(OR4_93_Y));
    OR4 OR4_744 (.A(\R_DATA_TEMPR44[13] ), .B(\R_DATA_TEMPR45[13] ), 
        .C(\R_DATA_TEMPR46[13] ), .D(\R_DATA_TEMPR47[13] ), .Y(
        OR4_744_Y));
    OR4 OR4_616 (.A(\R_DATA_TEMPR36[16] ), .B(\R_DATA_TEMPR37[16] ), 
        .C(\R_DATA_TEMPR38[16] ), .D(\R_DATA_TEMPR39[16] ), .Y(
        OR4_616_Y));
    OR4 OR4_309 (.A(\R_DATA_TEMPR36[34] ), .B(\R_DATA_TEMPR37[34] ), 
        .C(\R_DATA_TEMPR38[34] ), .D(\R_DATA_TEMPR39[34] ), .Y(
        OR4_309_Y));
    OR4 OR4_582 (.A(OR4_24_Y), .B(OR4_577_Y), .C(OR4_608_Y), .D(
        OR4_253_Y), .Y(OR4_582_Y));
    OR4 OR4_24 (.A(\R_DATA_TEMPR48[38] ), .B(\R_DATA_TEMPR49[38] ), .C(
        \R_DATA_TEMPR50[38] ), .D(\R_DATA_TEMPR51[38] ), .Y(OR4_24_Y));
    OR4 OR4_8 (.A(\R_DATA_TEMPR40[38] ), .B(\R_DATA_TEMPR41[38] ), .C(
        \R_DATA_TEMPR42[38] ), .D(\R_DATA_TEMPR43[38] ), .Y(OR4_8_Y));
    OR4 OR4_379 (.A(\R_DATA_TEMPR52[6] ), .B(\R_DATA_TEMPR53[6] ), .C(
        \R_DATA_TEMPR54[6] ), .D(\R_DATA_TEMPR55[6] ), .Y(OR4_379_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[7]  (.A(CFG3_13_Y), .B(CFG2_0_Y)
        , .Y(\BLKY2[7] ));
    OR4 OR4_250 (.A(\R_DATA_TEMPR48[20] ), .B(\R_DATA_TEMPR49[20] ), 
        .C(\R_DATA_TEMPR50[20] ), .D(\R_DATA_TEMPR51[20] ), .Y(
        OR4_250_Y));
    OR4 OR4_557 (.A(\R_DATA_TEMPR20[37] ), .B(\R_DATA_TEMPR21[37] ), 
        .C(\R_DATA_TEMPR22[37] ), .D(\R_DATA_TEMPR23[37] ), .Y(
        OR4_557_Y));
    OR4 OR4_334 (.A(OR4_350_Y), .B(OR4_227_Y), .C(OR4_76_Y), .D(
        OR4_405_Y), .Y(OR4_334_Y));
    OR4 OR4_791 (.A(\R_DATA_TEMPR8[30] ), .B(\R_DATA_TEMPR9[30] ), .C(
        \R_DATA_TEMPR10[30] ), .D(\R_DATA_TEMPR11[30] ), .Y(OR4_791_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R58C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%58%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R58C0 (
        .A_DOUT({\R_DATA_TEMPR58[39] , \R_DATA_TEMPR58[38] , 
        \R_DATA_TEMPR58[37] , \R_DATA_TEMPR58[36] , 
        \R_DATA_TEMPR58[35] , \R_DATA_TEMPR58[34] , 
        \R_DATA_TEMPR58[33] , \R_DATA_TEMPR58[32] , 
        \R_DATA_TEMPR58[31] , \R_DATA_TEMPR58[30] , 
        \R_DATA_TEMPR58[29] , \R_DATA_TEMPR58[28] , 
        \R_DATA_TEMPR58[27] , \R_DATA_TEMPR58[26] , 
        \R_DATA_TEMPR58[25] , \R_DATA_TEMPR58[24] , 
        \R_DATA_TEMPR58[23] , \R_DATA_TEMPR58[22] , 
        \R_DATA_TEMPR58[21] , \R_DATA_TEMPR58[20] }), .B_DOUT({
        \R_DATA_TEMPR58[19] , \R_DATA_TEMPR58[18] , 
        \R_DATA_TEMPR58[17] , \R_DATA_TEMPR58[16] , 
        \R_DATA_TEMPR58[15] , \R_DATA_TEMPR58[14] , 
        \R_DATA_TEMPR58[13] , \R_DATA_TEMPR58[12] , 
        \R_DATA_TEMPR58[11] , \R_DATA_TEMPR58[10] , 
        \R_DATA_TEMPR58[9] , \R_DATA_TEMPR58[8] , \R_DATA_TEMPR58[7] , 
        \R_DATA_TEMPR58[6] , \R_DATA_TEMPR58[5] , \R_DATA_TEMPR58[4] , 
        \R_DATA_TEMPR58[3] , \R_DATA_TEMPR58[2] , \R_DATA_TEMPR58[1] , 
        \R_DATA_TEMPR58[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[58][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[14] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[14] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_131 (.A(\R_DATA_TEMPR0[33] ), .B(\R_DATA_TEMPR1[33] ), .C(
        \R_DATA_TEMPR2[33] ), .D(\R_DATA_TEMPR3[33] ), .Y(OR4_131_Y));
    OR4 OR4_584 (.A(\R_DATA_TEMPR60[6] ), .B(\R_DATA_TEMPR61[6] ), .C(
        \R_DATA_TEMPR62[6] ), .D(\R_DATA_TEMPR63[6] ), .Y(OR4_584_Y));
    OR4 OR4_659 (.A(\R_DATA_TEMPR52[7] ), .B(\R_DATA_TEMPR53[7] ), .C(
        \R_DATA_TEMPR54[7] ), .D(\R_DATA_TEMPR55[7] ), .Y(OR4_659_Y));
    OR4 OR4_596 (.A(\R_DATA_TEMPR32[24] ), .B(\R_DATA_TEMPR33[24] ), 
        .C(\R_DATA_TEMPR34[24] ), .D(\R_DATA_TEMPR35[24] ), .Y(
        OR4_596_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[8]  (.A(CFG3_7_Y), .B(CFG2_3_Y), 
        .Y(\BLKX2[8] ));
    OR4 \OR4_R_DATA[39]  (.A(OR4_442_Y), .B(OR4_273_Y), .C(OR4_210_Y), 
        .D(OR4_60_Y), .Y(R_DATA[39]));
    OR4 OR4_256 (.A(\R_DATA_TEMPR12[25] ), .B(\R_DATA_TEMPR13[25] ), 
        .C(\R_DATA_TEMPR14[25] ), .D(\R_DATA_TEMPR15[25] ), .Y(
        OR4_256_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R37C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%37%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R37C0 (
        .A_DOUT({\R_DATA_TEMPR37[39] , \R_DATA_TEMPR37[38] , 
        \R_DATA_TEMPR37[37] , \R_DATA_TEMPR37[36] , 
        \R_DATA_TEMPR37[35] , \R_DATA_TEMPR37[34] , 
        \R_DATA_TEMPR37[33] , \R_DATA_TEMPR37[32] , 
        \R_DATA_TEMPR37[31] , \R_DATA_TEMPR37[30] , 
        \R_DATA_TEMPR37[29] , \R_DATA_TEMPR37[28] , 
        \R_DATA_TEMPR37[27] , \R_DATA_TEMPR37[26] , 
        \R_DATA_TEMPR37[25] , \R_DATA_TEMPR37[24] , 
        \R_DATA_TEMPR37[23] , \R_DATA_TEMPR37[22] , 
        \R_DATA_TEMPR37[21] , \R_DATA_TEMPR37[20] }), .B_DOUT({
        \R_DATA_TEMPR37[19] , \R_DATA_TEMPR37[18] , 
        \R_DATA_TEMPR37[17] , \R_DATA_TEMPR37[16] , 
        \R_DATA_TEMPR37[15] , \R_DATA_TEMPR37[14] , 
        \R_DATA_TEMPR37[13] , \R_DATA_TEMPR37[12] , 
        \R_DATA_TEMPR37[11] , \R_DATA_TEMPR37[10] , 
        \R_DATA_TEMPR37[9] , \R_DATA_TEMPR37[8] , \R_DATA_TEMPR37[7] , 
        \R_DATA_TEMPR37[6] , \R_DATA_TEMPR37[5] , \R_DATA_TEMPR37[4] , 
        \R_DATA_TEMPR37[3] , \R_DATA_TEMPR37[2] , \R_DATA_TEMPR37[1] , 
        \R_DATA_TEMPR37[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[37][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[9] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[9] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_75 (.A(\R_DATA_TEMPR56[24] ), .B(\R_DATA_TEMPR57[24] ), .C(
        \R_DATA_TEMPR58[24] ), .D(\R_DATA_TEMPR59[24] ), .Y(OR4_75_Y));
    OR4 OR4_431 (.A(\R_DATA_TEMPR8[8] ), .B(\R_DATA_TEMPR9[8] ), .C(
        \R_DATA_TEMPR10[8] ), .D(\R_DATA_TEMPR11[8] ), .Y(OR4_431_Y));
    OR4 OR4_91 (.A(\R_DATA_TEMPR36[10] ), .B(\R_DATA_TEMPR37[10] ), .C(
        \R_DATA_TEMPR38[10] ), .D(\R_DATA_TEMPR39[10] ), .Y(OR4_91_Y));
    CFG3 #( .INIT(8'h40) )  CFG3_2 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_2_Y));
    OR4 OR4_124 (.A(\R_DATA_TEMPR24[10] ), .B(\R_DATA_TEMPR25[10] ), 
        .C(\R_DATA_TEMPR26[10] ), .D(\R_DATA_TEMPR27[10] ), .Y(
        OR4_124_Y));
    OR4 OR4_438 (.A(\R_DATA_TEMPR48[36] ), .B(\R_DATA_TEMPR49[36] ), 
        .C(\R_DATA_TEMPR50[36] ), .D(\R_DATA_TEMPR51[36] ), .Y(
        OR4_438_Y));
    OR4 OR4_709 (.A(\R_DATA_TEMPR8[15] ), .B(\R_DATA_TEMPR9[15] ), .C(
        \R_DATA_TEMPR10[15] ), .D(\R_DATA_TEMPR11[15] ), .Y(OR4_709_Y));
    OR4 OR4_381 (.A(\R_DATA_TEMPR24[31] ), .B(\R_DATA_TEMPR25[31] ), 
        .C(\R_DATA_TEMPR26[31] ), .D(\R_DATA_TEMPR27[31] ), .Y(
        OR4_381_Y));
    OR4 OR4_654 (.A(OR4_726_Y), .B(OR4_48_Y), .C(OR4_140_Y), .D(
        OR4_777_Y), .Y(OR4_654_Y));
    OR4 OR4_779 (.A(\R_DATA_TEMPR24[28] ), .B(\R_DATA_TEMPR25[28] ), 
        .C(\R_DATA_TEMPR26[28] ), .D(\R_DATA_TEMPR27[28] ), .Y(
        OR4_779_Y));
    OR4 OR4_480 (.A(OR4_693_Y), .B(OR4_257_Y), .C(OR4_242_Y), .D(
        OR4_621_Y), .Y(OR4_480_Y));
    OR4 OR4_503 (.A(\R_DATA_TEMPR40[21] ), .B(\R_DATA_TEMPR41[21] ), 
        .C(\R_DATA_TEMPR42[21] ), .D(\R_DATA_TEMPR43[21] ), .Y(
        OR4_503_Y));
    OR4 OR4_314 (.A(\R_DATA_TEMPR28[4] ), .B(\R_DATA_TEMPR29[4] ), .C(
        \R_DATA_TEMPR30[4] ), .D(\R_DATA_TEMPR31[4] ), .Y(OR4_314_Y));
    OR4 OR4_721 (.A(\R_DATA_TEMPR56[2] ), .B(\R_DATA_TEMPR57[2] ), .C(
        \R_DATA_TEMPR58[2] ), .D(\R_DATA_TEMPR59[2] ), .Y(OR4_721_Y));
    OR4 OR4_43 (.A(\R_DATA_TEMPR48[18] ), .B(\R_DATA_TEMPR49[18] ), .C(
        \R_DATA_TEMPR50[18] ), .D(\R_DATA_TEMPR51[18] ), .Y(OR4_43_Y));
    OR4 OR4_573 (.A(OR4_723_Y), .B(OR4_394_Y), .C(OR4_559_Y), .D(
        OR4_162_Y), .Y(OR4_573_Y));
    OR4 OR4_539 (.A(\R_DATA_TEMPR4[38] ), .B(\R_DATA_TEMPR5[38] ), .C(
        \R_DATA_TEMPR6[38] ), .D(\R_DATA_TEMPR7[38] ), .Y(OR4_539_Y));
    CFG1 #( .INIT(2'h1) )  \INVBLKX0[0]  (.A(W_ADDR[9]), .Y(\BLKX0[0] )
        );
    OR4 OR4_111 (.A(\R_DATA_TEMPR20[26] ), .B(\R_DATA_TEMPR21[26] ), 
        .C(\R_DATA_TEMPR22[26] ), .D(\R_DATA_TEMPR23[26] ), .Y(
        OR4_111_Y));
    OR4 OR4_598 (.A(\R_DATA_TEMPR32[28] ), .B(\R_DATA_TEMPR33[28] ), 
        .C(\R_DATA_TEMPR34[28] ), .D(\R_DATA_TEMPR35[28] ), .Y(
        OR4_598_Y));
    CFG3 #( .INIT(8'h8) )  CFG3_1 (.A(R_ADDR[13]), .B(R_ADDR[12]), .C(
        R_ADDR[11]), .Y(CFG3_1_Y));
    OR4 OR4_59 (.A(\R_DATA_TEMPR16[23] ), .B(\R_DATA_TEMPR17[23] ), .C(
        \R_DATA_TEMPR18[23] ), .D(\R_DATA_TEMPR19[23] ), .Y(OR4_59_Y));
    OR4 OR4_530 (.A(\R_DATA_TEMPR4[23] ), .B(\R_DATA_TEMPR5[23] ), .C(
        \R_DATA_TEMPR6[23] ), .D(\R_DATA_TEMPR7[23] ), .Y(OR4_530_Y));
    OR4 OR4_263 (.A(\R_DATA_TEMPR60[11] ), .B(\R_DATA_TEMPR61[11] ), 
        .C(\R_DATA_TEMPR62[11] ), .D(\R_DATA_TEMPR63[11] ), .Y(
        OR4_263_Y));
    OR4 OR4_526 (.A(\R_DATA_TEMPR0[2] ), .B(\R_DATA_TEMPR1[2] ), .C(
        \R_DATA_TEMPR2[2] ), .D(\R_DATA_TEMPR3[2] ), .Y(OR4_526_Y));
    OR4 OR4_445 (.A(\R_DATA_TEMPR20[25] ), .B(\R_DATA_TEMPR21[25] ), 
        .C(\R_DATA_TEMPR22[25] ), .D(\R_DATA_TEMPR23[25] ), .Y(
        OR4_445_Y));
    OR4 OR4_411 (.A(\R_DATA_TEMPR24[5] ), .B(\R_DATA_TEMPR25[5] ), .C(
        \R_DATA_TEMPR26[5] ), .D(\R_DATA_TEMPR27[5] ), .Y(OR4_411_Y));
    CFG3 #( .INIT(8'h2) )  CFG3_11 (.A(R_ADDR[13]), .B(R_ADDR[12]), .C(
        R_ADDR[11]), .Y(CFG3_11_Y));
    OR4 OR4_496 (.A(\R_DATA_TEMPR56[30] ), .B(\R_DATA_TEMPR57[30] ), 
        .C(\R_DATA_TEMPR58[30] ), .D(\R_DATA_TEMPR59[30] ), .Y(
        OR4_496_Y));
    OR4 OR4_418 (.A(\R_DATA_TEMPR16[9] ), .B(\R_DATA_TEMPR17[9] ), .C(
        \R_DATA_TEMPR18[9] ), .D(\R_DATA_TEMPR19[9] ), .Y(OR4_418_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%13%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R13C0 (
        .A_DOUT({\R_DATA_TEMPR13[39] , \R_DATA_TEMPR13[38] , 
        \R_DATA_TEMPR13[37] , \R_DATA_TEMPR13[36] , 
        \R_DATA_TEMPR13[35] , \R_DATA_TEMPR13[34] , 
        \R_DATA_TEMPR13[33] , \R_DATA_TEMPR13[32] , 
        \R_DATA_TEMPR13[31] , \R_DATA_TEMPR13[30] , 
        \R_DATA_TEMPR13[29] , \R_DATA_TEMPR13[28] , 
        \R_DATA_TEMPR13[27] , \R_DATA_TEMPR13[26] , 
        \R_DATA_TEMPR13[25] , \R_DATA_TEMPR13[24] , 
        \R_DATA_TEMPR13[23] , \R_DATA_TEMPR13[22] , 
        \R_DATA_TEMPR13[21] , \R_DATA_TEMPR13[20] }), .B_DOUT({
        \R_DATA_TEMPR13[19] , \R_DATA_TEMPR13[18] , 
        \R_DATA_TEMPR13[17] , \R_DATA_TEMPR13[16] , 
        \R_DATA_TEMPR13[15] , \R_DATA_TEMPR13[14] , 
        \R_DATA_TEMPR13[13] , \R_DATA_TEMPR13[12] , 
        \R_DATA_TEMPR13[11] , \R_DATA_TEMPR13[10] , 
        \R_DATA_TEMPR13[9] , \R_DATA_TEMPR13[8] , \R_DATA_TEMPR13[7] , 
        \R_DATA_TEMPR13[6] , \R_DATA_TEMPR13[5] , \R_DATA_TEMPR13[4] , 
        \R_DATA_TEMPR13[3] , \R_DATA_TEMPR13[2] , \R_DATA_TEMPR13[1] , 
        \R_DATA_TEMPR13[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[3] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 \OR4_R_DATA[0]  (.A(OR4_660_Y), .B(OR4_749_Y), .C(OR4_501_Y), 
        .D(OR4_654_Y), .Y(R_DATA[0]));
    OR4 OR4_389 (.A(\R_DATA_TEMPR32[34] ), .B(\R_DATA_TEMPR33[34] ), 
        .C(\R_DATA_TEMPR34[34] ), .D(\R_DATA_TEMPR35[34] ), .Y(
        OR4_389_Y));
    OR4 OR4_392 (.A(OR4_538_Y), .B(OR4_659_Y), .C(OR4_746_Y), .D(
        OR4_740_Y), .Y(OR4_392_Y));
    OR4 OR4_19 (.A(\R_DATA_TEMPR8[24] ), .B(\R_DATA_TEMPR9[24] ), .C(
        \R_DATA_TEMPR10[24] ), .D(\R_DATA_TEMPR11[24] ), .Y(OR4_19_Y));
    OR4 OR4_41 (.A(\R_DATA_TEMPR48[14] ), .B(\R_DATA_TEMPR49[14] ), .C(
        \R_DATA_TEMPR50[14] ), .D(\R_DATA_TEMPR51[14] ), .Y(OR4_41_Y));
    OR4 OR4_333 (.A(\R_DATA_TEMPR56[33] ), .B(\R_DATA_TEMPR57[33] ), 
        .C(\R_DATA_TEMPR58[33] ), .D(\R_DATA_TEMPR59[33] ), .Y(
        OR4_333_Y));
    OR4 OR4_730 (.A(\R_DATA_TEMPR4[24] ), .B(\R_DATA_TEMPR5[24] ), .C(
        \R_DATA_TEMPR6[24] ), .D(\R_DATA_TEMPR7[24] ), .Y(OR4_730_Y));
    OR4 OR4_519 (.A(\R_DATA_TEMPR52[35] ), .B(\R_DATA_TEMPR53[35] ), 
        .C(\R_DATA_TEMPR54[35] ), .D(\R_DATA_TEMPR55[35] ), .Y(
        OR4_519_Y));
    OR4 OR4_668 (.A(\R_DATA_TEMPR20[1] ), .B(\R_DATA_TEMPR21[1] ), .C(
        \R_DATA_TEMPR22[1] ), .D(\R_DATA_TEMPR23[1] ), .Y(OR4_668_Y));
    OR4 OR4_510 (.A(\R_DATA_TEMPR60[8] ), .B(\R_DATA_TEMPR61[8] ), .C(
        \R_DATA_TEMPR62[8] ), .D(\R_DATA_TEMPR63[8] ), .Y(OR4_510_Y));
    OR4 OR4_432 (.A(\R_DATA_TEMPR52[27] ), .B(\R_DATA_TEMPR53[27] ), 
        .C(\R_DATA_TEMPR54[27] ), .D(\R_DATA_TEMPR55[27] ), .Y(
        OR4_432_Y));
    OR4 OR4_444 (.A(\R_DATA_TEMPR16[17] ), .B(\R_DATA_TEMPR17[17] ), 
        .C(\R_DATA_TEMPR18[17] ), .D(\R_DATA_TEMPR19[17] ), .Y(
        OR4_444_Y));
    OR4 OR4_528 (.A(\R_DATA_TEMPR40[17] ), .B(\R_DATA_TEMPR41[17] ), 
        .C(\R_DATA_TEMPR42[17] ), .D(\R_DATA_TEMPR43[17] ), .Y(
        OR4_528_Y));
    OR4 OR4_52 (.A(\R_DATA_TEMPR4[35] ), .B(\R_DATA_TEMPR5[35] ), .C(
        \R_DATA_TEMPR6[35] ), .D(\R_DATA_TEMPR7[35] ), .Y(OR4_52_Y));
    OR4 OR4_662 (.A(\R_DATA_TEMPR28[11] ), .B(\R_DATA_TEMPR29[11] ), 
        .C(\R_DATA_TEMPR30[11] ), .D(\R_DATA_TEMPR31[11] ), .Y(
        OR4_662_Y));
    OR4 OR4_439 (.A(\R_DATA_TEMPR56[16] ), .B(\R_DATA_TEMPR57[16] ), 
        .C(\R_DATA_TEMPR58[16] ), .D(\R_DATA_TEMPR59[16] ), .Y(
        OR4_439_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R40C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%40%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R40C0 (
        .A_DOUT({\R_DATA_TEMPR40[39] , \R_DATA_TEMPR40[38] , 
        \R_DATA_TEMPR40[37] , \R_DATA_TEMPR40[36] , 
        \R_DATA_TEMPR40[35] , \R_DATA_TEMPR40[34] , 
        \R_DATA_TEMPR40[33] , \R_DATA_TEMPR40[32] , 
        \R_DATA_TEMPR40[31] , \R_DATA_TEMPR40[30] , 
        \R_DATA_TEMPR40[29] , \R_DATA_TEMPR40[28] , 
        \R_DATA_TEMPR40[27] , \R_DATA_TEMPR40[26] , 
        \R_DATA_TEMPR40[25] , \R_DATA_TEMPR40[24] , 
        \R_DATA_TEMPR40[23] , \R_DATA_TEMPR40[22] , 
        \R_DATA_TEMPR40[21] , \R_DATA_TEMPR40[20] }), .B_DOUT({
        \R_DATA_TEMPR40[19] , \R_DATA_TEMPR40[18] , 
        \R_DATA_TEMPR40[17] , \R_DATA_TEMPR40[16] , 
        \R_DATA_TEMPR40[15] , \R_DATA_TEMPR40[14] , 
        \R_DATA_TEMPR40[13] , \R_DATA_TEMPR40[12] , 
        \R_DATA_TEMPR40[11] , \R_DATA_TEMPR40[10] , 
        \R_DATA_TEMPR40[9] , \R_DATA_TEMPR40[8] , \R_DATA_TEMPR40[7] , 
        \R_DATA_TEMPR40[6] , \R_DATA_TEMPR40[5] , \R_DATA_TEMPR40[4] , 
        \R_DATA_TEMPR40[3] , \R_DATA_TEMPR40[2] , \R_DATA_TEMPR40[1] , 
        \R_DATA_TEMPR40[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[40][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[10] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[10] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_346 (.A(OR4_679_Y), .B(OR4_1_Y), .C(OR4_95_Y), .D(
        OR4_176_Y), .Y(OR4_346_Y));
    OR4 OR4_136 (.A(\R_DATA_TEMPR44[7] ), .B(\R_DATA_TEMPR45[7] ), .C(
        \R_DATA_TEMPR46[7] ), .D(\R_DATA_TEMPR47[7] ), .Y(OR4_136_Y));
    CFG1 #( .INIT(2'h1) )  \INVBLKX1[0]  (.A(W_ADDR[10]), .Y(
        \BLKX1[0] ));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R49C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%49%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R49C0 (
        .A_DOUT({\R_DATA_TEMPR49[39] , \R_DATA_TEMPR49[38] , 
        \R_DATA_TEMPR49[37] , \R_DATA_TEMPR49[36] , 
        \R_DATA_TEMPR49[35] , \R_DATA_TEMPR49[34] , 
        \R_DATA_TEMPR49[33] , \R_DATA_TEMPR49[32] , 
        \R_DATA_TEMPR49[31] , \R_DATA_TEMPR49[30] , 
        \R_DATA_TEMPR49[29] , \R_DATA_TEMPR49[28] , 
        \R_DATA_TEMPR49[27] , \R_DATA_TEMPR49[26] , 
        \R_DATA_TEMPR49[25] , \R_DATA_TEMPR49[24] , 
        \R_DATA_TEMPR49[23] , \R_DATA_TEMPR49[22] , 
        \R_DATA_TEMPR49[21] , \R_DATA_TEMPR49[20] }), .B_DOUT({
        \R_DATA_TEMPR49[19] , \R_DATA_TEMPR49[18] , 
        \R_DATA_TEMPR49[17] , \R_DATA_TEMPR49[16] , 
        \R_DATA_TEMPR49[15] , \R_DATA_TEMPR49[14] , 
        \R_DATA_TEMPR49[13] , \R_DATA_TEMPR49[12] , 
        \R_DATA_TEMPR49[11] , \R_DATA_TEMPR49[10] , 
        \R_DATA_TEMPR49[9] , \R_DATA_TEMPR49[8] , \R_DATA_TEMPR49[7] , 
        \R_DATA_TEMPR49[6] , \R_DATA_TEMPR49[5] , \R_DATA_TEMPR49[4] , 
        \R_DATA_TEMPR49[3] , \R_DATA_TEMPR49[2] , \R_DATA_TEMPR49[1] , 
        \R_DATA_TEMPR49[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[49][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[12] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[12] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_426 (.A(OR4_714_Y), .B(OR4_38_Y), .C(OR4_125_Y), .D(
        OR4_770_Y), .Y(OR4_426_Y));
    OR4 OR4_203 (.A(\R_DATA_TEMPR36[30] ), .B(\R_DATA_TEMPR37[30] ), 
        .C(\R_DATA_TEMPR38[30] ), .D(\R_DATA_TEMPR39[30] ), .Y(
        OR4_203_Y));
    OR4 OR4_290 (.A(\R_DATA_TEMPR32[9] ), .B(\R_DATA_TEMPR33[9] ), .C(
        \R_DATA_TEMPR34[9] ), .D(\R_DATA_TEMPR35[9] ), .Y(OR4_290_Y));
    OR4 OR4_597 (.A(\R_DATA_TEMPR28[36] ), .B(\R_DATA_TEMPR29[36] ), 
        .C(\R_DATA_TEMPR30[36] ), .D(\R_DATA_TEMPR31[36] ), .Y(
        OR4_597_Y));
    OR4 OR4_789 (.A(\R_DATA_TEMPR60[5] ), .B(\R_DATA_TEMPR61[5] ), .C(
        \R_DATA_TEMPR62[5] ), .D(\R_DATA_TEMPR63[5] ), .Y(OR4_789_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R46C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%46%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R46C0 (
        .A_DOUT({\R_DATA_TEMPR46[39] , \R_DATA_TEMPR46[38] , 
        \R_DATA_TEMPR46[37] , \R_DATA_TEMPR46[36] , 
        \R_DATA_TEMPR46[35] , \R_DATA_TEMPR46[34] , 
        \R_DATA_TEMPR46[33] , \R_DATA_TEMPR46[32] , 
        \R_DATA_TEMPR46[31] , \R_DATA_TEMPR46[30] , 
        \R_DATA_TEMPR46[29] , \R_DATA_TEMPR46[28] , 
        \R_DATA_TEMPR46[27] , \R_DATA_TEMPR46[26] , 
        \R_DATA_TEMPR46[25] , \R_DATA_TEMPR46[24] , 
        \R_DATA_TEMPR46[23] , \R_DATA_TEMPR46[22] , 
        \R_DATA_TEMPR46[21] , \R_DATA_TEMPR46[20] }), .B_DOUT({
        \R_DATA_TEMPR46[19] , \R_DATA_TEMPR46[18] , 
        \R_DATA_TEMPR46[17] , \R_DATA_TEMPR46[16] , 
        \R_DATA_TEMPR46[15] , \R_DATA_TEMPR46[14] , 
        \R_DATA_TEMPR46[13] , \R_DATA_TEMPR46[12] , 
        \R_DATA_TEMPR46[11] , \R_DATA_TEMPR46[10] , 
        \R_DATA_TEMPR46[9] , \R_DATA_TEMPR46[8] , \R_DATA_TEMPR46[7] , 
        \R_DATA_TEMPR46[6] , \R_DATA_TEMPR46[5] , \R_DATA_TEMPR46[4] , 
        \R_DATA_TEMPR46[3] , \R_DATA_TEMPR46[2] , \R_DATA_TEMPR46[1] , 
        \R_DATA_TEMPR46[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[46][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[11] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[11] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_338 (.A(\R_DATA_TEMPR16[30] ), .B(\R_DATA_TEMPR17[30] ), 
        .C(\R_DATA_TEMPR18[30] ), .D(\R_DATA_TEMPR19[30] ), .Y(
        OR4_338_Y));
    OR4 OR4_273 (.A(OR4_617_Y), .B(OR4_649_Y), .C(OR4_638_Y), .D(
        OR4_479_Y), .Y(OR4_273_Y));
    OR4 OR4_313 (.A(\R_DATA_TEMPR44[31] ), .B(\R_DATA_TEMPR45[31] ), 
        .C(\R_DATA_TEMPR46[31] ), .D(\R_DATA_TEMPR47[31] ), .Y(
        OR4_313_Y));
    OR4 OR4_322 (.A(\R_DATA_TEMPR8[29] ), .B(\R_DATA_TEMPR9[29] ), .C(
        \R_DATA_TEMPR10[29] ), .D(\R_DATA_TEMPR11[29] ), .Y(OR4_322_Y));
    OR4 OR4_710 (.A(OR4_642_Y), .B(OR4_115_Y), .C(OR4_503_Y), .D(
        OR4_637_Y), .Y(OR4_710_Y));
    OR4 OR4_699 (.A(\R_DATA_TEMPR56[22] ), .B(\R_DATA_TEMPR57[22] ), 
        .C(\R_DATA_TEMPR58[22] ), .D(\R_DATA_TEMPR59[22] ), .Y(
        OR4_699_Y));
    OR4 OR4_12 (.A(\R_DATA_TEMPR36[25] ), .B(\R_DATA_TEMPR37[25] ), .C(
        \R_DATA_TEMPR38[25] ), .D(\R_DATA_TEMPR39[25] ), .Y(OR4_12_Y));
    CFG3 #( .INIT(8'h40) )  CFG3_12 (.A(R_ADDR[13]), .B(R_ADDR[12]), 
        .C(R_ADDR[11]), .Y(CFG3_12_Y));
    OR4 OR4_583 (.A(\R_DATA_TEMPR8[7] ), .B(\R_DATA_TEMPR9[7] ), .C(
        \R_DATA_TEMPR10[7] ), .D(\R_DATA_TEMPR11[7] ), .Y(OR4_583_Y));
    OR4 OR4_412 (.A(\R_DATA_TEMPR28[25] ), .B(\R_DATA_TEMPR29[25] ), 
        .C(\R_DATA_TEMPR30[25] ), .D(\R_DATA_TEMPR31[25] ), .Y(
        OR4_412_Y));
    OR4 OR4_296 (.A(\R_DATA_TEMPR44[4] ), .B(\R_DATA_TEMPR45[4] ), .C(
        \R_DATA_TEMPR46[4] ), .D(\R_DATA_TEMPR47[4] ), .Y(OR4_296_Y));
    OR4 OR4_419 (.A(\R_DATA_TEMPR60[2] ), .B(\R_DATA_TEMPR61[2] ), .C(
        \R_DATA_TEMPR62[2] ), .D(\R_DATA_TEMPR63[2] ), .Y(OR4_419_Y));
    OR4 OR4_251 (.A(\R_DATA_TEMPR4[2] ), .B(\R_DATA_TEMPR5[2] ), .C(
        \R_DATA_TEMPR6[2] ), .D(\R_DATA_TEMPR7[2] ), .Y(OR4_251_Y));
    OR4 OR4_79 (.A(\R_DATA_TEMPR44[32] ), .B(\R_DATA_TEMPR45[32] ), .C(
        \R_DATA_TEMPR46[32] ), .D(\R_DATA_TEMPR47[32] ), .Y(OR4_79_Y));
    OR4 OR4_139 (.A(\R_DATA_TEMPR20[10] ), .B(\R_DATA_TEMPR21[10] ), 
        .C(\R_DATA_TEMPR22[10] ), .D(\R_DATA_TEMPR23[10] ), .Y(
        OR4_139_Y));
    OR4 OR4_116 (.A(\R_DATA_TEMPR56[21] ), .B(\R_DATA_TEMPR57[21] ), 
        .C(\R_DATA_TEMPR58[21] ), .D(\R_DATA_TEMPR59[21] ), .Y(
        OR4_116_Y));
    OR4 OR4_608 (.A(\R_DATA_TEMPR56[38] ), .B(\R_DATA_TEMPR57[38] ), 
        .C(\R_DATA_TEMPR58[38] ), .D(\R_DATA_TEMPR59[38] ), .Y(
        OR4_608_Y));
    OR4 OR4_144 (.A(OR4_701_Y), .B(OR4_539_Y), .C(OR4_404_Y), .D(
        OR4_443_Y), .Y(OR4_144_Y));
    OR4 OR4_694 (.A(OR4_449_Y), .B(OR4_292_Y), .C(OR4_151_Y), .D(
        OR4_190_Y), .Y(OR4_694_Y));
    OR4 OR4_678 (.A(\R_DATA_TEMPR4[17] ), .B(\R_DATA_TEMPR5[17] ), .C(
        \R_DATA_TEMPR6[17] ), .D(\R_DATA_TEMPR7[17] ), .Y(OR4_678_Y));
    OR4 OR4_602 (.A(\R_DATA_TEMPR32[37] ), .B(\R_DATA_TEMPR33[37] ), 
        .C(\R_DATA_TEMPR34[37] ), .D(\R_DATA_TEMPR35[37] ), .Y(
        OR4_602_Y));
    OR4 \OR4_R_DATA[32]  (.A(OR4_762_Y), .B(OR4_735_Y), .C(OR4_627_Y), 
        .D(OR4_279_Y), .Y(R_DATA[32]));
    OR4 OR4_552 (.A(OR4_444_Y), .B(OR4_458_Y), .C(OR4_448_Y), .D(
        OR4_29_Y), .Y(OR4_552_Y));
    OR4 OR4_220 (.A(\R_DATA_TEMPR16[7] ), .B(\R_DATA_TEMPR17[7] ), .C(
        \R_DATA_TEMPR18[7] ), .D(\R_DATA_TEMPR19[7] ), .Y(OR4_220_Y));
    OR4 OR4_672 (.A(\R_DATA_TEMPR60[35] ), .B(\R_DATA_TEMPR61[35] ), 
        .C(\R_DATA_TEMPR62[35] ), .D(\R_DATA_TEMPR63[35] ), .Y(
        OR4_672_Y));
    OR4 OR4_527 (.A(\R_DATA_TEMPR0[20] ), .B(\R_DATA_TEMPR1[20] ), .C(
        \R_DATA_TEMPR2[20] ), .D(\R_DATA_TEMPR3[20] ), .Y(OR4_527_Y));
    OR4 OR4_318 (.A(\R_DATA_TEMPR56[19] ), .B(\R_DATA_TEMPR57[19] ), 
        .C(\R_DATA_TEMPR58[19] ), .D(\R_DATA_TEMPR59[19] ), .Y(
        OR4_318_Y));
    OR4 OR4_741 (.A(\R_DATA_TEMPR24[7] ), .B(\R_DATA_TEMPR25[7] ), .C(
        \R_DATA_TEMPR26[7] ), .D(\R_DATA_TEMPR27[7] ), .Y(OR4_741_Y));
    OR4 \OR4_R_DATA[3]  (.A(OR4_194_Y), .B(OR4_415_Y), .C(OR4_354_Y), 
        .D(OR4_413_Y), .Y(R_DATA[3]));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%18%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R18C0 (
        .A_DOUT({\R_DATA_TEMPR18[39] , \R_DATA_TEMPR18[38] , 
        \R_DATA_TEMPR18[37] , \R_DATA_TEMPR18[36] , 
        \R_DATA_TEMPR18[35] , \R_DATA_TEMPR18[34] , 
        \R_DATA_TEMPR18[33] , \R_DATA_TEMPR18[32] , 
        \R_DATA_TEMPR18[31] , \R_DATA_TEMPR18[30] , 
        \R_DATA_TEMPR18[29] , \R_DATA_TEMPR18[28] , 
        \R_DATA_TEMPR18[27] , \R_DATA_TEMPR18[26] , 
        \R_DATA_TEMPR18[25] , \R_DATA_TEMPR18[24] , 
        \R_DATA_TEMPR18[23] , \R_DATA_TEMPR18[22] , 
        \R_DATA_TEMPR18[21] , \R_DATA_TEMPR18[20] }), .B_DOUT({
        \R_DATA_TEMPR18[19] , \R_DATA_TEMPR18[18] , 
        \R_DATA_TEMPR18[17] , \R_DATA_TEMPR18[16] , 
        \R_DATA_TEMPR18[15] , \R_DATA_TEMPR18[14] , 
        \R_DATA_TEMPR18[13] , \R_DATA_TEMPR18[12] , 
        \R_DATA_TEMPR18[11] , \R_DATA_TEMPR18[10] , 
        \R_DATA_TEMPR18[9] , \R_DATA_TEMPR18[8] , \R_DATA_TEMPR18[7] , 
        \R_DATA_TEMPR18[6] , \R_DATA_TEMPR18[5] , \R_DATA_TEMPR18[4] , 
        \R_DATA_TEMPR18[3] , \R_DATA_TEMPR18[2] , \R_DATA_TEMPR18[1] , 
        \R_DATA_TEMPR18[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[4] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[4] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_666 (.A(\R_DATA_TEMPR32[12] ), .B(\R_DATA_TEMPR33[12] ), 
        .C(\R_DATA_TEMPR34[12] ), .D(\R_DATA_TEMPR35[12] ), .Y(
        OR4_666_Y));
    OR4 OR4_629 (.A(\R_DATA_TEMPR16[24] ), .B(\R_DATA_TEMPR17[24] ), 
        .C(\R_DATA_TEMPR18[24] ), .D(\R_DATA_TEMPR19[24] ), .Y(
        OR4_629_Y));
    OR4 OR4_554 (.A(OR4_219_Y), .B(OR4_58_Y), .C(OR4_49_Y), .D(
        OR4_440_Y), .Y(OR4_554_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R63C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%63%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R63C0 (
        .A_DOUT({\R_DATA_TEMPR63[39] , \R_DATA_TEMPR63[38] , 
        \R_DATA_TEMPR63[37] , \R_DATA_TEMPR63[36] , 
        \R_DATA_TEMPR63[35] , \R_DATA_TEMPR63[34] , 
        \R_DATA_TEMPR63[33] , \R_DATA_TEMPR63[32] , 
        \R_DATA_TEMPR63[31] , \R_DATA_TEMPR63[30] , 
        \R_DATA_TEMPR63[29] , \R_DATA_TEMPR63[28] , 
        \R_DATA_TEMPR63[27] , \R_DATA_TEMPR63[26] , 
        \R_DATA_TEMPR63[25] , \R_DATA_TEMPR63[24] , 
        \R_DATA_TEMPR63[23] , \R_DATA_TEMPR63[22] , 
        \R_DATA_TEMPR63[21] , \R_DATA_TEMPR63[20] }), .B_DOUT({
        \R_DATA_TEMPR63[19] , \R_DATA_TEMPR63[18] , 
        \R_DATA_TEMPR63[17] , \R_DATA_TEMPR63[16] , 
        \R_DATA_TEMPR63[15] , \R_DATA_TEMPR63[14] , 
        \R_DATA_TEMPR63[13] , \R_DATA_TEMPR63[12] , 
        \R_DATA_TEMPR63[11] , \R_DATA_TEMPR63[10] , 
        \R_DATA_TEMPR63[9] , \R_DATA_TEMPR63[8] , \R_DATA_TEMPR63[7] , 
        \R_DATA_TEMPR63[6] , \R_DATA_TEMPR63[5] , \R_DATA_TEMPR63[4] , 
        \R_DATA_TEMPR63[3] , \R_DATA_TEMPR63[2] , \R_DATA_TEMPR63[1] , 
        \R_DATA_TEMPR63[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[63][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[15] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[15] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_546 (.A(\R_DATA_TEMPR24[37] ), .B(\R_DATA_TEMPR25[37] ), 
        .C(\R_DATA_TEMPR26[37] ), .D(\R_DATA_TEMPR27[37] ), .Y(
        OR4_546_Y));
    OR4 OR4_226 (.A(\R_DATA_TEMPR52[24] ), .B(\R_DATA_TEMPR53[24] ), 
        .C(\R_DATA_TEMPR54[24] ), .D(\R_DATA_TEMPR55[24] ), .Y(
        OR4_226_Y));
    OR4 OR4_119 (.A(\R_DATA_TEMPR20[9] ), .B(\R_DATA_TEMPR21[9] ), .C(
        \R_DATA_TEMPR22[9] ), .D(\R_DATA_TEMPR23[9] ), .Y(OR4_119_Y));
    OR4 OR4_72 (.A(\R_DATA_TEMPR36[28] ), .B(\R_DATA_TEMPR37[28] ), .C(
        \R_DATA_TEMPR38[28] ), .D(\R_DATA_TEMPR39[28] ), .Y(OR4_72_Y));
    OR4 OR4_735 (.A(OR4_399_Y), .B(OR4_169_Y), .C(OR4_158_Y), .D(
        OR4_799_Y), .Y(OR4_735_Y));
    OR4 OR4_637 (.A(\R_DATA_TEMPR44[21] ), .B(\R_DATA_TEMPR45[21] ), 
        .C(\R_DATA_TEMPR46[21] ), .D(\R_DATA_TEMPR47[21] ), .Y(
        OR4_637_Y));
    OR4 OR4_736 (.A(OR4_120_Y), .B(OR4_111_Y), .C(OR4_383_Y), .D(
        OR4_83_Y), .Y(OR4_736_Y));
    OR4 OR4_624 (.A(\R_DATA_TEMPR52[31] ), .B(\R_DATA_TEMPR53[31] ), 
        .C(\R_DATA_TEMPR54[31] ), .D(\R_DATA_TEMPR55[31] ), .Y(
        OR4_624_Y));
    OR4 OR4_351 (.A(\R_DATA_TEMPR20[34] ), .B(\R_DATA_TEMPR21[34] ), 
        .C(\R_DATA_TEMPR22[34] ), .D(\R_DATA_TEMPR23[34] ), .Y(
        OR4_351_Y));
    OR4 \OR4_R_DATA[33]  (.A(OR4_675_Y), .B(OR4_462_Y), .C(OR4_436_Y), 
        .D(OR4_407_Y), .Y(R_DATA[33]));
    OR4 \OR4_R_DATA[25]  (.A(OR4_633_Y), .B(OR4_216_Y), .C(OR4_524_Y), 
        .D(OR4_301_Y), .Y(R_DATA[25]));
    OR4 OR4_450 (.A(\R_DATA_TEMPR20[2] ), .B(\R_DATA_TEMPR21[2] ), .C(
        \R_DATA_TEMPR22[2] ), .D(\R_DATA_TEMPR23[2] ), .Y(OR4_450_Y));
    OR4 OR4_283 (.A(\R_DATA_TEMPR0[11] ), .B(\R_DATA_TEMPR1[11] ), .C(
        \R_DATA_TEMPR2[11] ), .D(\R_DATA_TEMPR3[11] ), .Y(OR4_283_Y));
    OR4 OR4_96 (.A(\R_DATA_TEMPR12[39] ), .B(\R_DATA_TEMPR13[39] ), .C(
        \R_DATA_TEMPR14[39] ), .D(\R_DATA_TEMPR15[39] ), .Y(OR4_96_Y));
    OR4 OR4_548 (.A(\R_DATA_TEMPR48[33] ), .B(\R_DATA_TEMPR49[33] ), 
        .C(\R_DATA_TEMPR50[33] ), .D(\R_DATA_TEMPR51[33] ), .Y(
        OR4_548_Y));
    OR4 OR4_54 (.A(\R_DATA_TEMPR16[4] ), .B(\R_DATA_TEMPR17[4] ), .C(
        \R_DATA_TEMPR18[4] ), .D(\R_DATA_TEMPR19[4] ), .Y(OR4_54_Y));
    OR4 OR4_3 (.A(\R_DATA_TEMPR52[11] ), .B(\R_DATA_TEMPR53[11] ), .C(
        \R_DATA_TEMPR54[11] ), .D(\R_DATA_TEMPR55[11] ), .Y(OR4_3_Y));
    OR4 OR4_364 (.A(\R_DATA_TEMPR28[0] ), .B(\R_DATA_TEMPR29[0] ), .C(
        \R_DATA_TEMPR30[0] ), .D(\R_DATA_TEMPR31[0] ), .Y(OR4_364_Y));
    OR4 OR4_606 (.A(\R_DATA_TEMPR4[30] ), .B(\R_DATA_TEMPR5[30] ), .C(
        \R_DATA_TEMPR6[30] ), .D(\R_DATA_TEMPR7[30] ), .Y(OR4_606_Y));
    OR4 OR4_715 (.A(\R_DATA_TEMPR20[27] ), .B(\R_DATA_TEMPR21[27] ), 
        .C(\R_DATA_TEMPR22[27] ), .D(\R_DATA_TEMPR23[27] ), .Y(
        OR4_715_Y));
    OR4 OR4_617 (.A(\R_DATA_TEMPR16[39] ), .B(\R_DATA_TEMPR17[39] ), 
        .C(\R_DATA_TEMPR18[39] ), .D(\R_DATA_TEMPR19[39] ), .Y(
        OR4_617_Y));
    OR4 OR4_161 (.A(\R_DATA_TEMPR44[30] ), .B(\R_DATA_TEMPR45[30] ), 
        .C(\R_DATA_TEMPR46[30] ), .D(\R_DATA_TEMPR47[30] ), .Y(
        OR4_161_Y));
    OR4 OR4_446 (.A(OR4_666_Y), .B(OR4_16_Y), .C(OR4_128_Y), .D(
        OR4_39_Y), .Y(OR4_446_Y));
    OR4 OR4_716 (.A(\R_DATA_TEMPR40[0] ), .B(\R_DATA_TEMPR41[0] ), .C(
        \R_DATA_TEMPR42[0] ), .D(\R_DATA_TEMPR43[0] ), .Y(OR4_716_Y));
    OR4 OR4_676 (.A(\R_DATA_TEMPR40[27] ), .B(\R_DATA_TEMPR41[27] ), 
        .C(\R_DATA_TEMPR42[27] ), .D(\R_DATA_TEMPR43[27] ), .Y(
        OR4_676_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[6]  (.A(CFG3_1_Y), .B(CFG2_0_Y), 
        .Y(\BLKY2[6] ));
    OR4 OR4_237 (.A(\R_DATA_TEMPR16[18] ), .B(\R_DATA_TEMPR17[18] ), 
        .C(\R_DATA_TEMPR18[18] ), .D(\R_DATA_TEMPR19[18] ), .Y(
        OR4_237_Y));
    OR4 OR4_688 (.A(\R_DATA_TEMPR28[6] ), .B(\R_DATA_TEMPR29[6] ), .C(
        \R_DATA_TEMPR30[6] ), .D(\R_DATA_TEMPR31[6] ), .Y(OR4_688_Y));
    OR4 OR4_137 (.A(\R_DATA_TEMPR60[37] ), .B(\R_DATA_TEMPR61[37] ), 
        .C(\R_DATA_TEMPR62[37] ), .D(\R_DATA_TEMPR63[37] ), .Y(
        OR4_137_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%2%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R2C0 (.A_DOUT({
        \R_DATA_TEMPR2[39] , \R_DATA_TEMPR2[38] , \R_DATA_TEMPR2[37] , 
        \R_DATA_TEMPR2[36] , \R_DATA_TEMPR2[35] , \R_DATA_TEMPR2[34] , 
        \R_DATA_TEMPR2[33] , \R_DATA_TEMPR2[32] , \R_DATA_TEMPR2[31] , 
        \R_DATA_TEMPR2[30] , \R_DATA_TEMPR2[29] , \R_DATA_TEMPR2[28] , 
        \R_DATA_TEMPR2[27] , \R_DATA_TEMPR2[26] , \R_DATA_TEMPR2[25] , 
        \R_DATA_TEMPR2[24] , \R_DATA_TEMPR2[23] , \R_DATA_TEMPR2[22] , 
        \R_DATA_TEMPR2[21] , \R_DATA_TEMPR2[20] }), .B_DOUT({
        \R_DATA_TEMPR2[19] , \R_DATA_TEMPR2[18] , \R_DATA_TEMPR2[17] , 
        \R_DATA_TEMPR2[16] , \R_DATA_TEMPR2[15] , \R_DATA_TEMPR2[14] , 
        \R_DATA_TEMPR2[13] , \R_DATA_TEMPR2[12] , \R_DATA_TEMPR2[11] , 
        \R_DATA_TEMPR2[10] , \R_DATA_TEMPR2[9] , \R_DATA_TEMPR2[8] , 
        \R_DATA_TEMPR2[7] , \R_DATA_TEMPR2[6] , \R_DATA_TEMPR2[5] , 
        \R_DATA_TEMPR2[4] , \R_DATA_TEMPR2[3] , \R_DATA_TEMPR2[2] , 
        \R_DATA_TEMPR2[1] , \R_DATA_TEMPR2[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[2][0] ), .A_ADDR({
        R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[0] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_682 (.A(\R_DATA_TEMPR24[8] ), .B(\R_DATA_TEMPR25[8] ), .C(
        \R_DATA_TEMPR26[8] ), .D(\R_DATA_TEMPR27[8] ), .Y(OR4_682_Y));
    OR4 OR4_342 (.A(\R_DATA_TEMPR4[21] ), .B(\R_DATA_TEMPR5[21] ), .C(
        \R_DATA_TEMPR6[21] ), .D(\R_DATA_TEMPR7[21] ), .Y(OR4_342_Y));
    OR4 OR4_359 (.A(\R_DATA_TEMPR40[20] ), .B(\R_DATA_TEMPR41[20] ), 
        .C(\R_DATA_TEMPR42[20] ), .D(\R_DATA_TEMPR43[20] ), .Y(
        OR4_359_Y));
    OR4 OR4_461 (.A(OR4_150_Y), .B(OR4_293_Y), .C(OR4_284_Y), .D(
        OR4_109_Y), .Y(OR4_461_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[11]  (.A(CFG3_2_Y), .B(CFG2_3_Y)
        , .Y(\BLKX2[11] ));
    OR4 OR4_14 (.A(\R_DATA_TEMPR0[34] ), .B(\R_DATA_TEMPR1[34] ), .C(
        \R_DATA_TEMPR2[34] ), .D(\R_DATA_TEMPR3[34] ), .Y(OR4_14_Y));
    OR4 OR4_468 (.A(\R_DATA_TEMPR60[39] ), .B(\R_DATA_TEMPR61[39] ), 
        .C(\R_DATA_TEMPR62[39] ), .D(\R_DATA_TEMPR63[39] ), .Y(
        OR4_468_Y));
    OR4 OR4_733 (.A(OR4_625_Y), .B(OR4_557_Y), .C(OR4_546_Y), .D(
        OR4_388_Y), .Y(OR4_733_Y));
    OR4 OR4_291 (.A(\R_DATA_TEMPR48[25] ), .B(\R_DATA_TEMPR49[25] ), 
        .C(\R_DATA_TEMPR50[25] ), .D(\R_DATA_TEMPR51[25] ), .Y(
        OR4_291_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R33C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%33%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R33C0 (
        .A_DOUT({\R_DATA_TEMPR33[39] , \R_DATA_TEMPR33[38] , 
        \R_DATA_TEMPR33[37] , \R_DATA_TEMPR33[36] , 
        \R_DATA_TEMPR33[35] , \R_DATA_TEMPR33[34] , 
        \R_DATA_TEMPR33[33] , \R_DATA_TEMPR33[32] , 
        \R_DATA_TEMPR33[31] , \R_DATA_TEMPR33[30] , 
        \R_DATA_TEMPR33[29] , \R_DATA_TEMPR33[28] , 
        \R_DATA_TEMPR33[27] , \R_DATA_TEMPR33[26] , 
        \R_DATA_TEMPR33[25] , \R_DATA_TEMPR33[24] , 
        \R_DATA_TEMPR33[23] , \R_DATA_TEMPR33[22] , 
        \R_DATA_TEMPR33[21] , \R_DATA_TEMPR33[20] }), .B_DOUT({
        \R_DATA_TEMPR33[19] , \R_DATA_TEMPR33[18] , 
        \R_DATA_TEMPR33[17] , \R_DATA_TEMPR33[16] , 
        \R_DATA_TEMPR33[15] , \R_DATA_TEMPR33[14] , 
        \R_DATA_TEMPR33[13] , \R_DATA_TEMPR33[12] , 
        \R_DATA_TEMPR33[11] , \R_DATA_TEMPR33[10] , 
        \R_DATA_TEMPR33[9] , \R_DATA_TEMPR33[8] , \R_DATA_TEMPR33[7] , 
        \R_DATA_TEMPR33[6] , \R_DATA_TEMPR33[5] , \R_DATA_TEMPR33[4] , 
        \R_DATA_TEMPR33[3] , \R_DATA_TEMPR33[2] , \R_DATA_TEMPR33[1] , 
        \R_DATA_TEMPR33[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[33][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[8] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[8] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_234 (.A(\R_DATA_TEMPR60[24] ), .B(\R_DATA_TEMPR61[24] ), 
        .C(\R_DATA_TEMPR62[24] ), .D(\R_DATA_TEMPR63[24] ), .Y(
        OR4_234_Y));
    OR4 OR4_90 (.A(\R_DATA_TEMPR8[35] ), .B(\R_DATA_TEMPR9[35] ), .C(
        \R_DATA_TEMPR10[35] ), .D(\R_DATA_TEMPR11[35] ), .Y(OR4_90_Y));
    OR4 OR4_46 (.A(\R_DATA_TEMPR60[12] ), .B(\R_DATA_TEMPR61[12] ), .C(
        \R_DATA_TEMPR62[12] ), .D(\R_DATA_TEMPR63[12] ), .Y(OR4_46_Y));
    OR4 OR4_569 (.A(\R_DATA_TEMPR32[13] ), .B(\R_DATA_TEMPR33[13] ), 
        .C(\R_DATA_TEMPR34[13] ), .D(\R_DATA_TEMPR35[13] ), .Y(
        OR4_569_Y));
    OR4 OR4_97 (.A(\R_DATA_TEMPR8[4] ), .B(\R_DATA_TEMPR9[4] ), .C(
        \R_DATA_TEMPR10[4] ), .D(\R_DATA_TEMPR11[4] ), .Y(OR4_97_Y));
    OR4 \OR4_R_DATA[6]  (.A(OR4_187_Y), .B(OR4_565_Y), .C(OR4_30_Y), 
        .D(OR4_134_Y), .Y(R_DATA[6]));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R42C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%42%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R42C0 (
        .A_DOUT({\R_DATA_TEMPR42[39] , \R_DATA_TEMPR42[38] , 
        \R_DATA_TEMPR42[37] , \R_DATA_TEMPR42[36] , 
        \R_DATA_TEMPR42[35] , \R_DATA_TEMPR42[34] , 
        \R_DATA_TEMPR42[33] , \R_DATA_TEMPR42[32] , 
        \R_DATA_TEMPR42[31] , \R_DATA_TEMPR42[30] , 
        \R_DATA_TEMPR42[29] , \R_DATA_TEMPR42[28] , 
        \R_DATA_TEMPR42[27] , \R_DATA_TEMPR42[26] , 
        \R_DATA_TEMPR42[25] , \R_DATA_TEMPR42[24] , 
        \R_DATA_TEMPR42[23] , \R_DATA_TEMPR42[22] , 
        \R_DATA_TEMPR42[21] , \R_DATA_TEMPR42[20] }), .B_DOUT({
        \R_DATA_TEMPR42[19] , \R_DATA_TEMPR42[18] , 
        \R_DATA_TEMPR42[17] , \R_DATA_TEMPR42[16] , 
        \R_DATA_TEMPR42[15] , \R_DATA_TEMPR42[14] , 
        \R_DATA_TEMPR42[13] , \R_DATA_TEMPR42[12] , 
        \R_DATA_TEMPR42[11] , \R_DATA_TEMPR42[10] , 
        \R_DATA_TEMPR42[9] , \R_DATA_TEMPR42[8] , \R_DATA_TEMPR42[7] , 
        \R_DATA_TEMPR42[6] , \R_DATA_TEMPR42[5] , \R_DATA_TEMPR42[4] , 
        \R_DATA_TEMPR42[3] , \R_DATA_TEMPR42[2] , \R_DATA_TEMPR42[1] , 
        \R_DATA_TEMPR42[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[42][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[10] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[10] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], 
        W_DATA[16], W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], 
        W_DATA[11], W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], 
        W_DATA[6], W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], 
        W_DATA[1], W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], 
        WBYTE_EN[0]}), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        VCC, GND, VCC}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_592 (.A(\R_DATA_TEMPR0[10] ), .B(\R_DATA_TEMPR1[10] ), .C(
        \R_DATA_TEMPR2[10] ), .D(\R_DATA_TEMPR3[10] ), .Y(OR4_592_Y));
    OR4 OR4_63 (.A(\R_DATA_TEMPR52[39] ), .B(\R_DATA_TEMPR53[39] ), .C(
        \R_DATA_TEMPR54[39] ), .D(\R_DATA_TEMPR55[39] ), .Y(OR4_63_Y));
    OR4 OR4_560 (.A(\R_DATA_TEMPR8[16] ), .B(\R_DATA_TEMPR9[16] ), .C(
        \R_DATA_TEMPR10[16] ), .D(\R_DATA_TEMPR11[16] ), .Y(OR4_560_Y));
    OR4 OR4_217 (.A(OR4_59_Y), .B(OR4_241_Y), .C(OR4_497_Y), .D(
        OR4_206_Y), .Y(OR4_217_Y));
    OR4 OR4_240 (.A(\R_DATA_TEMPR0[17] ), .B(\R_DATA_TEMPR1[17] ), .C(
        \R_DATA_TEMPR2[17] ), .D(\R_DATA_TEMPR3[17] ), .Y(OR4_240_Y));
    OR4 OR4_304 (.A(\R_DATA_TEMPR52[9] ), .B(\R_DATA_TEMPR53[9] ), .C(
        \R_DATA_TEMPR54[9] ), .D(\R_DATA_TEMPR55[9] ), .Y(OR4_304_Y));
    OR4 OR4_117 (.A(OR4_758_Y), .B(OR4_639_Y), .C(OR4_491_Y), .D(
        OR4_551_Y), .Y(OR4_117_Y));
    OR4 OR4_547 (.A(\R_DATA_TEMPR20[21] ), .B(\R_DATA_TEMPR21[21] ), 
        .C(\R_DATA_TEMPR22[21] ), .D(\R_DATA_TEMPR23[21] ), .Y(
        OR4_547_Y));
    OR4 OR4_335 (.A(\R_DATA_TEMPR44[0] ), .B(\R_DATA_TEMPR45[0] ), .C(
        \R_DATA_TEMPR46[0] ), .D(\R_DATA_TEMPR47[0] ), .Y(OR4_335_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[3]  (.A(CFG3_12_Y), .B(CFG2_0_Y)
        , .Y(\BLKY2[3] ));
    OR4 OR4_374 (.A(\R_DATA_TEMPR16[27] ), .B(\R_DATA_TEMPR17[27] ), 
        .C(\R_DATA_TEMPR18[27] ), .D(\R_DATA_TEMPR19[27] ), .Y(
        OR4_374_Y));
    OR4 \OR4_R_DATA[1]  (.A(OR4_652_Y), .B(OR4_743_Y), .C(OR4_533_Y), 
        .D(OR4_426_Y), .Y(R_DATA[1]));
    OR4 OR4_101 (.A(OR4_259_Y), .B(OR4_702_Y), .C(OR4_447_Y), .D(
        OR4_174_Y), .Y(OR4_101_Y));
    OR4 OR4_759 (.A(OR4_121_Y), .B(OR4_147_Y), .C(OR4_411_Y), .D(
        OR4_634_Y), .Y(OR4_759_Y));
    OR4 OR4_649 (.A(\R_DATA_TEMPR20[39] ), .B(\R_DATA_TEMPR21[39] ), 
        .C(\R_DATA_TEMPR22[39] ), .D(\R_DATA_TEMPR23[39] ), .Y(
        OR4_649_Y));
    OR4 OR4_594 (.A(\R_DATA_TEMPR4[31] ), .B(\R_DATA_TEMPR5[31] ), .C(
        \R_DATA_TEMPR6[31] ), .D(\R_DATA_TEMPR7[31] ), .Y(OR4_594_Y));
    OR4 OR4_171 (.A(\R_DATA_TEMPR28[7] ), .B(\R_DATA_TEMPR29[7] ), .C(
        \R_DATA_TEMPR30[7] ), .D(\R_DATA_TEMPR31[7] ), .Y(OR4_171_Y));
    OR4 OR4_713 (.A(\R_DATA_TEMPR12[19] ), .B(\R_DATA_TEMPR13[19] ), 
        .C(\R_DATA_TEMPR14[19] ), .D(\R_DATA_TEMPR15[19] ), .Y(
        OR4_713_Y));
    OR4 OR4_553 (.A(\R_DATA_TEMPR28[15] ), .B(\R_DATA_TEMPR29[15] ), 
        .C(\R_DATA_TEMPR30[15] ), .D(\R_DATA_TEMPR31[15] ), .Y(
        OR4_553_Y));
    OR4 OR4_214 (.A(\R_DATA_TEMPR40[10] ), .B(\R_DATA_TEMPR41[10] ), 
        .C(\R_DATA_TEMPR42[10] ), .D(\R_DATA_TEMPR43[10] ), .Y(
        OR4_214_Y));
    OR4 OR4_246 (.A(\R_DATA_TEMPR36[11] ), .B(\R_DATA_TEMPR37[11] ), 
        .C(\R_DATA_TEMPR38[11] ), .D(\R_DATA_TEMPR39[11] ), .Y(
        OR4_246_Y));
    OR4 OR4_221 (.A(\R_DATA_TEMPR56[36] ), .B(\R_DATA_TEMPR57[36] ), 
        .C(\R_DATA_TEMPR58[36] ), .D(\R_DATA_TEMPR59[36] ), .Y(
        OR4_221_Y));
    OR4 OR4_401 (.A(OR4_43_Y), .B(OR4_764_Y), .C(OR4_27_Y), .D(
        OR4_143_Y), .Y(OR4_401_Y));
    OR4 OR4_74 (.A(OR4_393_Y), .B(OR4_52_Y), .C(OR4_90_Y), .D(
        OR4_498_Y), .Y(OR4_74_Y));
    OR4 OR4_408 (.A(\R_DATA_TEMPR8[11] ), .B(\R_DATA_TEMPR9[11] ), .C(
        \R_DATA_TEMPR10[11] ), .D(\R_DATA_TEMPR11[11] ), .Y(OR4_408_Y));
    OR4 OR4_732 (.A(\R_DATA_TEMPR48[10] ), .B(\R_DATA_TEMPR49[10] ), 
        .C(\R_DATA_TEMPR50[10] ), .D(\R_DATA_TEMPR51[10] ), .Y(
        OR4_732_Y));
    OR4 OR4_471 (.A(\R_DATA_TEMPR12[21] ), .B(\R_DATA_TEMPR13[21] ), 
        .C(\R_DATA_TEMPR14[21] ), .D(\R_DATA_TEMPR15[21] ), .Y(
        OR4_471_Y));
    OR4 OR4_363 (.A(OR4_788_Y), .B(OR4_698_Y), .C(OR4_754_Y), .D(
        OR4_563_Y), .Y(OR4_363_Y));
    OR4 OR4_760 (.A(OR4_522_Y), .B(OR4_352_Y), .C(OR4_222_Y), .D(
        OR4_269_Y), .Y(OR4_760_Y));
    OR4 OR4_478 (.A(\R_DATA_TEMPR16[1] ), .B(\R_DATA_TEMPR17[1] ), .C(
        \R_DATA_TEMPR18[1] ), .D(\R_DATA_TEMPR19[1] ), .Y(OR4_478_Y));
    OR4 OR4_391 (.A(\R_DATA_TEMPR32[38] ), .B(\R_DATA_TEMPR33[38] ), 
        .C(\R_DATA_TEMPR34[38] ), .D(\R_DATA_TEMPR35[38] ), .Y(
        OR4_391_Y));
    OR4 OR4_644 (.A(\R_DATA_TEMPR48[32] ), .B(\R_DATA_TEMPR49[32] ), 
        .C(\R_DATA_TEMPR50[32] ), .D(\R_DATA_TEMPR51[32] ), .Y(
        OR4_644_Y));
    OR4 OR4_61 (.A(\R_DATA_TEMPR60[34] ), .B(\R_DATA_TEMPR61[34] ), .C(
        \R_DATA_TEMPR62[34] ), .D(\R_DATA_TEMPR63[34] ), .Y(OR4_61_Y));
    OR4 OR4_462 (.A(OR4_321_Y), .B(OR4_69_Y), .C(OR4_57_Y), .D(
        OR4_711_Y), .Y(OR4_462_Y));
    OR4 OR4_635 (.A(\R_DATA_TEMPR0[14] ), .B(\R_DATA_TEMPR1[14] ), .C(
        \R_DATA_TEMPR2[14] ), .D(\R_DATA_TEMPR3[14] ), .Y(OR4_635_Y));
    OR4 OR4_522 (.A(\R_DATA_TEMPR0[18] ), .B(\R_DATA_TEMPR1[18] ), .C(
        \R_DATA_TEMPR2[18] ), .D(\R_DATA_TEMPR3[18] ), .Y(OR4_522_Y));
    OR4 OR4_686 (.A(OR4_336_Y), .B(OR4_267_Y), .C(OR4_318_Y), .D(
        OR4_367_Y), .Y(OR4_686_Y));
    OR4 OR4_315 (.A(\R_DATA_TEMPR48[39] ), .B(\R_DATA_TEMPR49[39] ), 
        .C(\R_DATA_TEMPR50[39] ), .D(\R_DATA_TEMPR51[39] ), .Y(
        OR4_315_Y));
    OR4 OR4_469 (.A(\R_DATA_TEMPR56[6] ), .B(\R_DATA_TEMPR57[6] ), .C(
        \R_DATA_TEMPR58[6] ), .D(\R_DATA_TEMPR59[6] ), .Y(OR4_469_Y));
    OR4 OR4_490 (.A(\R_DATA_TEMPR40[2] ), .B(\R_DATA_TEMPR41[2] ), .C(
        \R_DATA_TEMPR42[2] ), .D(\R_DATA_TEMPR43[2] ), .Y(OR4_490_Y));
    OR4 OR4_40 (.A(\R_DATA_TEMPR4[19] ), .B(\R_DATA_TEMPR5[19] ), .C(
        \R_DATA_TEMPR6[19] ), .D(\R_DATA_TEMPR7[19] ), .Y(OR4_40_Y));
    OR4 OR4_509 (.A(OR4_648_Y), .B(OR4_794_Y), .C(OR4_525_Y), .D(
        OR4_136_Y), .Y(OR4_509_Y));
    OR4 OR4_166 (.A(\R_DATA_TEMPR48[22] ), .B(\R_DATA_TEMPR49[22] ), 
        .C(\R_DATA_TEMPR50[22] ), .D(\R_DATA_TEMPR51[22] ), .Y(
        OR4_166_Y));
    OR4 OR4_500 (.A(\R_DATA_TEMPR48[2] ), .B(\R_DATA_TEMPR49[2] ), .C(
        \R_DATA_TEMPR50[2] ), .D(\R_DATA_TEMPR51[2] ), .Y(OR4_500_Y));
    OR4 OR4_47 (.A(\R_DATA_TEMPR32[18] ), .B(\R_DATA_TEMPR33[18] ), .C(
        \R_DATA_TEMPR34[18] ), .D(\R_DATA_TEMPR35[18] ), .Y(OR4_47_Y));
    OR4 OR4_579 (.A(\R_DATA_TEMPR44[9] ), .B(\R_DATA_TEMPR45[9] ), .C(
        \R_DATA_TEMPR46[9] ), .D(\R_DATA_TEMPR47[9] ), .Y(OR4_579_Y));
    OR4 OR4_570 (.A(\R_DATA_TEMPR32[8] ), .B(\R_DATA_TEMPR33[8] ), .C(
        \R_DATA_TEMPR34[8] ), .D(\R_DATA_TEMPR35[8] ), .Y(OR4_570_Y));
    OR4 OR4_524 (.A(OR4_536_Y), .B(OR4_12_Y), .C(OR4_400_Y), .D(
        OR4_529_Y), .Y(OR4_524_Y));
    OR4 \OR4_R_DATA[28]  (.A(OR4_694_Y), .B(OR4_587_Y), .C(OR4_229_Y), 
        .D(OR4_334_Y), .Y(R_DATA[28]));
    OR4 OR4_368 (.A(\R_DATA_TEMPR28[20] ), .B(\R_DATA_TEMPR29[20] ), 
        .C(\R_DATA_TEMPR30[20] ), .D(\R_DATA_TEMPR31[20] ), .Y(
        OR4_368_Y));
    OR4 OR4_712 (.A(OR4_55_Y), .B(OR4_624_Y), .C(OR4_651_Y), .D(
        OR4_355_Y), .Y(OR4_712_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R38C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%38%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R38C0 (
        .A_DOUT({\R_DATA_TEMPR38[39] , \R_DATA_TEMPR38[38] , 
        \R_DATA_TEMPR38[37] , \R_DATA_TEMPR38[36] , 
        \R_DATA_TEMPR38[35] , \R_DATA_TEMPR38[34] , 
        \R_DATA_TEMPR38[33] , \R_DATA_TEMPR38[32] , 
        \R_DATA_TEMPR38[31] , \R_DATA_TEMPR38[30] , 
        \R_DATA_TEMPR38[29] , \R_DATA_TEMPR38[28] , 
        \R_DATA_TEMPR38[27] , \R_DATA_TEMPR38[26] , 
        \R_DATA_TEMPR38[25] , \R_DATA_TEMPR38[24] , 
        \R_DATA_TEMPR38[23] , \R_DATA_TEMPR38[22] , 
        \R_DATA_TEMPR38[21] , \R_DATA_TEMPR38[20] }), .B_DOUT({
        \R_DATA_TEMPR38[19] , \R_DATA_TEMPR38[18] , 
        \R_DATA_TEMPR38[17] , \R_DATA_TEMPR38[16] , 
        \R_DATA_TEMPR38[15] , \R_DATA_TEMPR38[14] , 
        \R_DATA_TEMPR38[13] , \R_DATA_TEMPR38[12] , 
        \R_DATA_TEMPR38[11] , \R_DATA_TEMPR38[10] , 
        \R_DATA_TEMPR38[9] , \R_DATA_TEMPR38[8] , \R_DATA_TEMPR38[7] , 
        \R_DATA_TEMPR38[6] , \R_DATA_TEMPR38[5] , \R_DATA_TEMPR38[4] , 
        \R_DATA_TEMPR38[3] , \R_DATA_TEMPR38[2] , \R_DATA_TEMPR38[1] , 
        \R_DATA_TEMPR38[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[38][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[9] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[9] , W_ADDR[10], \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_630 (.A(\R_DATA_TEMPR52[2] ), .B(\R_DATA_TEMPR53[2] ), .C(
        \R_DATA_TEMPR54[2] ), .D(\R_DATA_TEMPR55[2] ), .Y(OR4_630_Y));
    RAM1K20 #( .MEMORYFILE("PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C0.mem")
        , .RAMINDEX("PF_SRAM_AHB_C0%32768-32768%40-40%POWER%24%0%TWO-PORT%hex/miv-rv32i-systick-blinky.hex%ECC_EN-0")
         )  PF_SRAM_AHB_C0_PF_TPSRAM_AHB_AXI_0_PF_TPSRAM_R24C0 (
        .A_DOUT({\R_DATA_TEMPR24[39] , \R_DATA_TEMPR24[38] , 
        \R_DATA_TEMPR24[37] , \R_DATA_TEMPR24[36] , 
        \R_DATA_TEMPR24[35] , \R_DATA_TEMPR24[34] , 
        \R_DATA_TEMPR24[33] , \R_DATA_TEMPR24[32] , 
        \R_DATA_TEMPR24[31] , \R_DATA_TEMPR24[30] , 
        \R_DATA_TEMPR24[29] , \R_DATA_TEMPR24[28] , 
        \R_DATA_TEMPR24[27] , \R_DATA_TEMPR24[26] , 
        \R_DATA_TEMPR24[25] , \R_DATA_TEMPR24[24] , 
        \R_DATA_TEMPR24[23] , \R_DATA_TEMPR24[22] , 
        \R_DATA_TEMPR24[21] , \R_DATA_TEMPR24[20] }), .B_DOUT({
        \R_DATA_TEMPR24[19] , \R_DATA_TEMPR24[18] , 
        \R_DATA_TEMPR24[17] , \R_DATA_TEMPR24[16] , 
        \R_DATA_TEMPR24[15] , \R_DATA_TEMPR24[14] , 
        \R_DATA_TEMPR24[13] , \R_DATA_TEMPR24[12] , 
        \R_DATA_TEMPR24[11] , \R_DATA_TEMPR24[10] , 
        \R_DATA_TEMPR24[9] , \R_DATA_TEMPR24[8] , \R_DATA_TEMPR24[7] , 
        \R_DATA_TEMPR24[6] , \R_DATA_TEMPR24[5] , \R_DATA_TEMPR24[4] , 
        \R_DATA_TEMPR24[3] , \R_DATA_TEMPR24[2] , \R_DATA_TEMPR24[1] , 
        \R_DATA_TEMPR24[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[24][0] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({W_DATA[39], W_DATA[38], W_DATA[37], W_DATA[36], 
        W_DATA[35], W_DATA[34], W_DATA[33], W_DATA[32], W_DATA[31], 
        W_DATA[30], W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], 
        W_DATA[25], W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], 
        W_DATA[20]}), .A_REN(VCC), .A_WEN({WBYTE_EN[3], WBYTE_EN[2]}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[6] , \BLKX1[0] , \BLKX0[0] }), .B_CLK(
        CLK), .B_DIN({W_DATA[19], W_DATA[18], W_DATA[17], W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({WBYTE_EN[1], WBYTE_EN[0]}), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_98 (.A(\R_DATA_TEMPR56[39] ), .B(\R_DATA_TEMPR57[39] ), .C(
        \R_DATA_TEMPR58[39] ), .D(\R_DATA_TEMPR59[39] ), .Y(OR4_98_Y));
    OR4 OR4_321 (.A(\R_DATA_TEMPR16[33] ), .B(\R_DATA_TEMPR17[33] ), 
        .C(\R_DATA_TEMPR18[33] ), .D(\R_DATA_TEMPR19[33] ), .Y(
        OR4_321_Y));
    OR4 OR4_615 (.A(\R_DATA_TEMPR4[27] ), .B(\R_DATA_TEMPR5[27] ), .C(
        \R_DATA_TEMPR6[27] ), .D(\R_DATA_TEMPR7[27] ), .Y(OR4_615_Y));
    OR4 OR4_337 (.A(\R_DATA_TEMPR32[19] ), .B(\R_DATA_TEMPR33[19] ), 
        .C(\R_DATA_TEMPR34[19] ), .D(\R_DATA_TEMPR35[19] ), .Y(
        OR4_337_Y));
    OR4 OR4_130 (.A(\R_DATA_TEMPR36[4] ), .B(\R_DATA_TEMPR37[4] ), .C(
        \R_DATA_TEMPR38[4] ), .D(\R_DATA_TEMPR39[4] ), .Y(OR4_130_Y));
    OR4 OR4_169 (.A(\R_DATA_TEMPR20[32] ), .B(\R_DATA_TEMPR21[32] ), 
        .C(\R_DATA_TEMPR22[32] ), .D(\R_DATA_TEMPR23[32] ), .Y(
        OR4_169_Y));
    OR4 OR4_303 (.A(OR4_570_Y), .B(OR4_724_Y), .C(OR4_455_Y), .D(
        OR4_64_Y), .Y(OR4_303_Y));
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule
